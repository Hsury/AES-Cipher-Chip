
module aes_encipher_block ( clk, reset_n, next, keylen, round, round_key, 
        sboxw, new_sboxw, block, new_block, ready );
  output [3:0] round;
  input [127:0] round_key;
  output [31:0] sboxw;
  input [31:0] new_sboxw;
  input [127:0] block;
  output [127:0] new_block;
  input clk, reset_n, next, keylen;
  output ready;
  wire   enc_ctrl_we, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1222, n1223,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n256, n1221, n1224, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463;
  wire   [1:0] sword_ctr_reg;
  wire   [2:0] enc_ctrl_reg;

  DFFSX1 ready_reg_reg ( .D(n1361), .CK(clk), .SN(n1382), .Q(ready) );
  DFFRX1 \block_w1_reg_reg[23]  ( .D(n1272), .CK(clk), .RN(n1382), .Q(
        new_block[87]), .QN(n91) );
  DFFRX1 \block_w2_reg_reg[23]  ( .D(n1304), .CK(clk), .RN(n1381), .Q(
        new_block[55]), .QN(n59) );
  DFFRX1 \block_w0_reg_reg[22]  ( .D(n1242), .CK(clk), .RN(n1382), .Q(
        new_block[118]), .QN(n124) );
  DFFRX1 \block_w0_reg_reg[23]  ( .D(n1241), .CK(clk), .RN(n1384), .Q(
        new_block[119]), .QN(n123) );
  DFFRX1 \block_w3_reg_reg[22]  ( .D(n1337), .CK(clk), .RN(n1379), .Q(
        new_block[22]), .QN(n22) );
  DFFRX1 \block_w3_reg_reg[23]  ( .D(n1336), .CK(clk), .RN(n1381), .Q(
        new_block[23]), .QN(n21) );
  DFFRX1 \block_w1_reg_reg[31]  ( .D(n1264), .CK(clk), .RN(n1380), .Q(
        new_block[95]), .QN(n83) );
  DFFRX1 \block_w2_reg_reg[31]  ( .D(n1296), .CK(clk), .RN(n1380), .Q(
        new_block[63]), .QN(n51) );
  DFFRX1 \block_w0_reg_reg[31]  ( .D(n1233), .CK(clk), .RN(n1372), .Q(
        new_block[127]), .QN(n115) );
  DFFRX1 \block_w3_reg_reg[31]  ( .D(n1328), .CK(clk), .RN(n1381), .Q(
        new_block[31]), .QN(n13) );
  DFFRX1 \block_w1_reg_reg[22]  ( .D(n1273), .CK(clk), .RN(n1371), .Q(
        new_block[86]), .QN(n92) );
  DFFRX1 \block_w1_reg_reg[21]  ( .D(n1274), .CK(clk), .RN(n1384), .Q(
        new_block[85]), .QN(n93) );
  DFFRX1 \block_w2_reg_reg[22]  ( .D(n1305), .CK(clk), .RN(n1380), .Q(
        new_block[54]), .QN(n60) );
  DFFRX1 \block_w2_reg_reg[21]  ( .D(n1306), .CK(clk), .RN(n1381), .Q(
        new_block[53]), .QN(n61) );
  DFFRX1 \block_w0_reg_reg[21]  ( .D(n1243), .CK(clk), .RN(n1383), .Q(
        new_block[117]), .QN(n125) );
  DFFRX1 \block_w3_reg_reg[21]  ( .D(n1338), .CK(clk), .RN(n1383), .Q(
        new_block[21]), .QN(n23) );
  DFFRX1 \block_w1_reg_reg[29]  ( .D(n1266), .CK(clk), .RN(n1372), .Q(
        new_block[93]), .QN(n85) );
  DFFRX1 \block_w1_reg_reg[30]  ( .D(n1265), .CK(clk), .RN(n1371), .Q(
        new_block[94]), .QN(n84) );
  DFFRX1 \block_w2_reg_reg[30]  ( .D(n1297), .CK(clk), .RN(n1382), .Q(
        new_block[62]), .QN(n52) );
  DFFRX1 \block_w0_reg_reg[29]  ( .D(n1235), .CK(clk), .RN(n1372), .Q(
        new_block[125]), .QN(n117) );
  DFFRX1 \block_w0_reg_reg[30]  ( .D(n1234), .CK(clk), .RN(n1382), .Q(
        new_block[126]), .QN(n116) );
  DFFRX1 \block_w3_reg_reg[30]  ( .D(n1329), .CK(clk), .RN(n1371), .Q(
        new_block[30]), .QN(n14) );
  DFFRX1 \block_w3_reg_reg[29]  ( .D(n1330), .CK(clk), .RN(n1381), .Q(
        new_block[29]), .QN(n15) );
  DFFRX1 \round_ctr_reg_reg[0]  ( .D(n1365), .CK(clk), .RN(n1373), .Q(round[0]), .QN(n48) );
  DFFRX1 \block_w1_reg_reg[16]  ( .D(n1279), .CK(clk), .RN(n1383), .Q(
        new_block[80]), .QN(n98) );
  DFFRX1 \block_w1_reg_reg[17]  ( .D(n1278), .CK(clk), .RN(n1370), .Q(
        new_block[81]), .QN(n97) );
  DFFRX1 \block_w1_reg_reg[18]  ( .D(n1277), .CK(clk), .RN(n1383), .Q(
        new_block[82]), .QN(n96) );
  DFFRX1 \block_w1_reg_reg[19]  ( .D(n1276), .CK(clk), .RN(n1384), .Q(
        new_block[83]), .QN(n95) );
  DFFRX1 \block_w1_reg_reg[20]  ( .D(n1275), .CK(clk), .RN(n1370), .Q(
        new_block[84]), .QN(n94) );
  DFFRX1 \block_w2_reg_reg[17]  ( .D(n1310), .CK(clk), .RN(n1384), .Q(
        new_block[49]), .QN(n65) );
  DFFRX1 \block_w2_reg_reg[20]  ( .D(n1307), .CK(clk), .RN(n1370), .Q(
        new_block[52]), .QN(n62) );
  DFFRX1 \block_w0_reg_reg[20]  ( .D(n1244), .CK(clk), .RN(n1370), .Q(
        new_block[116]), .QN(n126) );
  DFFRX1 \block_w0_reg_reg[17]  ( .D(n1247), .CK(clk), .RN(n1383), .Q(
        new_block[113]), .QN(n129) );
  DFFRX1 \block_w3_reg_reg[20]  ( .D(n1339), .CK(clk), .RN(n1370), .Q(
        new_block[20]), .QN(n24) );
  DFFRX1 \block_w3_reg_reg[17]  ( .D(n1342), .CK(clk), .RN(n1382), .Q(
        new_block[17]), .QN(n27) );
  DFFRX1 \block_w2_reg_reg[16]  ( .D(n1311), .CK(clk), .RN(n1382), .Q(
        new_block[48]), .QN(n66) );
  DFFRX1 \block_w2_reg_reg[18]  ( .D(n1309), .CK(clk), .RN(n1381), .Q(
        new_block[50]), .QN(n64) );
  DFFRX1 \block_w2_reg_reg[19]  ( .D(n1308), .CK(clk), .RN(n1370), .Q(
        new_block[51]), .QN(n63) );
  DFFRX1 \block_w0_reg_reg[18]  ( .D(n1246), .CK(clk), .RN(n1384), .Q(
        new_block[114]), .QN(n128) );
  DFFRX1 \block_w0_reg_reg[19]  ( .D(n1245), .CK(clk), .RN(n1370), .Q(
        new_block[115]), .QN(n127) );
  DFFRX1 \block_w0_reg_reg[16]  ( .D(n1248), .CK(clk), .RN(n1378), .Q(
        new_block[112]), .QN(n130) );
  DFFRX1 \block_w3_reg_reg[18]  ( .D(n1341), .CK(clk), .RN(n1383), .Q(
        new_block[18]), .QN(n26) );
  DFFRX1 \block_w3_reg_reg[19]  ( .D(n1340), .CK(clk), .RN(n1370), .Q(
        new_block[19]), .QN(n25) );
  DFFRX1 \block_w3_reg_reg[16]  ( .D(n1343), .CK(clk), .RN(n1381), .Q(
        new_block[16]), .QN(n28) );
  DFFRX1 \block_w1_reg_reg[28]  ( .D(n1267), .CK(clk), .RN(n1380), .Q(
        new_block[92]), .QN(n86) );
  DFFRX1 \block_w2_reg_reg[25]  ( .D(n1302), .CK(clk), .RN(n1372), .Q(
        new_block[57]), .QN(n57) );
  DFFRX1 \block_w2_reg_reg[28]  ( .D(n1299), .CK(clk), .RN(n1381), .Q(
        new_block[60]), .QN(n54) );
  DFFRX1 \block_w2_reg_reg[29]  ( .D(n1298), .CK(clk), .RN(n1384), .Q(
        new_block[61]), .QN(n53) );
  DFFRX1 \block_w1_reg_reg[24]  ( .D(n1271), .CK(clk), .RN(n1380), .Q(
        new_block[88]), .QN(n90) );
  DFFRX1 \block_w1_reg_reg[25]  ( .D(n1270), .CK(clk), .RN(n1380), .Q(
        new_block[89]), .QN(n89) );
  DFFRX1 \block_w1_reg_reg[26]  ( .D(n1269), .CK(clk), .RN(n1380), .Q(
        new_block[90]), .QN(n88) );
  DFFRX1 \block_w1_reg_reg[27]  ( .D(n1268), .CK(clk), .RN(n1380), .Q(
        new_block[91]), .QN(n87) );
  DFFRX1 \block_w2_reg_reg[26]  ( .D(n1301), .CK(clk), .RN(n1372), .Q(
        new_block[58]), .QN(n56) );
  DFFRX1 \block_w2_reg_reg[27]  ( .D(n1300), .CK(clk), .RN(n1383), .Q(
        new_block[59]), .QN(n55) );
  DFFRX1 \block_w2_reg_reg[24]  ( .D(n1303), .CK(clk), .RN(n1382), .Q(
        new_block[56]), .QN(n58) );
  DFFRX1 \block_w0_reg_reg[26]  ( .D(n1238), .CK(clk), .RN(n1371), .Q(
        new_block[122]), .QN(n120) );
  DFFRX1 \block_w0_reg_reg[24]  ( .D(n1240), .CK(clk), .RN(n1372), .Q(
        new_block[120]), .QN(n122) );
  DFFRX1 \block_w0_reg_reg[25]  ( .D(n1239), .CK(clk), .RN(n1371), .Q(
        new_block[121]), .QN(n121) );
  DFFRX1 \block_w0_reg_reg[28]  ( .D(n1236), .CK(clk), .RN(n1372), .Q(
        new_block[124]), .QN(n118) );
  DFFRX1 \block_w3_reg_reg[26]  ( .D(n1333), .CK(clk), .RN(n1384), .Q(
        new_block[26]), .QN(n18) );
  DFFRX1 \block_w3_reg_reg[24]  ( .D(n1335), .CK(clk), .RN(n1371), .Q(
        new_block[24]), .QN(n20) );
  DFFRX1 \block_w3_reg_reg[25]  ( .D(n1334), .CK(clk), .RN(n1383), .Q(
        new_block[25]), .QN(n19) );
  DFFRX1 \block_w3_reg_reg[28]  ( .D(n1331), .CK(clk), .RN(n1370), .Q(
        new_block[28]), .QN(n16) );
  DFFRX1 \block_w0_reg_reg[27]  ( .D(n1237), .CK(clk), .RN(n1372), .Q(
        new_block[123]), .QN(n119) );
  DFFRX1 \block_w3_reg_reg[27]  ( .D(n1332), .CK(clk), .RN(n1370), .Q(
        new_block[27]), .QN(n17) );
  DFFRX1 \block_w1_reg_reg[7]  ( .D(n1288), .CK(clk), .RN(n1378), .Q(
        new_block[71]), .QN(n107) );
  DFFRX1 \block_w2_reg_reg[7]  ( .D(n1320), .CK(clk), .RN(n1378), .Q(
        new_block[39]), .QN(n75) );
  DFFRX1 \block_w0_reg_reg[6]  ( .D(n1258), .CK(clk), .RN(n1377), .Q(
        new_block[102]), .QN(n140) );
  DFFRX1 \block_w0_reg_reg[7]  ( .D(n1257), .CK(clk), .RN(n1377), .Q(
        new_block[103]), .QN(n139) );
  DFFRX1 \block_w3_reg_reg[6]  ( .D(n1353), .CK(clk), .RN(n1377), .Q(
        new_block[6]), .QN(n38) );
  DFFRX1 \block_w3_reg_reg[7]  ( .D(n1352), .CK(clk), .RN(n1377), .Q(
        new_block[7]), .QN(n37) );
  DFFRX1 \block_w1_reg_reg[6]  ( .D(n1289), .CK(clk), .RN(n1377), .Q(
        new_block[70]), .QN(n108) );
  DFFRX1 \block_w2_reg_reg[6]  ( .D(n1321), .CK(clk), .RN(n1377), .Q(
        new_block[38]), .QN(n76) );
  DFFRX1 \block_w3_reg_reg[4]  ( .D(n1355), .CK(clk), .RN(n1376), .Q(
        new_block[4]), .QN(n40) );
  DFFRX1 \block_w0_reg_reg[15]  ( .D(n1249), .CK(clk), .RN(n1377), .Q(
        new_block[111]), .QN(n131) );
  DFFRX1 \block_w3_reg_reg[15]  ( .D(n1344), .CK(clk), .RN(n1378), .Q(
        new_block[15]), .QN(n29) );
  DFFRX1 \block_w0_reg_reg[4]  ( .D(n1260), .CK(clk), .RN(n1376), .Q(
        new_block[100]), .QN(n142) );
  DFFRX1 \block_w1_reg_reg[4]  ( .D(n1291), .CK(clk), .RN(n1376), .Q(
        new_block[68]), .QN(n110) );
  DFFRX1 \block_w2_reg_reg[4]  ( .D(n1323), .CK(clk), .RN(n1376), .Q(
        new_block[36]), .QN(n78) );
  DFFRX1 \block_w1_reg_reg[15]  ( .D(n1280), .CK(clk), .RN(n1377), .Q(
        new_block[79]), .QN(n99) );
  DFFRX1 \block_w2_reg_reg[15]  ( .D(n1312), .CK(clk), .RN(n1378), .Q(
        new_block[47]), .QN(n67) );
  DFFRX1 \block_w1_reg_reg[1]  ( .D(n1294), .CK(clk), .RN(n1374), .Q(
        new_block[65]), .QN(n113) );
  DFFRX1 \block_w2_reg_reg[1]  ( .D(n1326), .CK(clk), .RN(n1374), .Q(
        new_block[33]), .QN(n81) );
  DFFRX1 \block_w1_reg_reg[0]  ( .D(n1295), .CK(clk), .RN(n1373), .Q(
        new_block[64]), .QN(n114) );
  DFFRX1 \block_w1_reg_reg[2]  ( .D(n1293), .CK(clk), .RN(n1375), .Q(
        new_block[66]), .QN(n112) );
  DFFRX1 \block_w1_reg_reg[3]  ( .D(n1292), .CK(clk), .RN(n1375), .Q(
        new_block[67]), .QN(n111) );
  DFFRX1 \block_w1_reg_reg[5]  ( .D(n1290), .CK(clk), .RN(n1376), .Q(
        new_block[69]), .QN(n109) );
  DFFRX1 \block_w2_reg_reg[5]  ( .D(n1322), .CK(clk), .RN(n1377), .Q(
        new_block[37]), .QN(n77) );
  DFFRX1 \block_w3_reg_reg[1]  ( .D(n1358), .CK(clk), .RN(n1374), .Q(
        new_block[1]), .QN(n43) );
  DFFRX1 \block_w3_reg_reg[5]  ( .D(n1354), .CK(clk), .RN(n1377), .Q(
        new_block[5]), .QN(n39) );
  DFFRX1 \block_w0_reg_reg[1]  ( .D(n1263), .CK(clk), .RN(n1374), .Q(
        new_block[97]), .QN(n145) );
  DFFRX1 \block_w0_reg_reg[2]  ( .D(n1262), .CK(clk), .RN(n1375), .Q(
        new_block[98]), .QN(n144) );
  DFFRX1 \block_w0_reg_reg[3]  ( .D(n1261), .CK(clk), .RN(n1375), .Q(
        new_block[99]), .QN(n143) );
  DFFRX1 \block_w0_reg_reg[5]  ( .D(n1259), .CK(clk), .RN(n1376), .Q(
        new_block[101]), .QN(n141) );
  DFFRX1 \block_w2_reg_reg[0]  ( .D(n1327), .CK(clk), .RN(n1374), .Q(
        new_block[32]), .QN(n82) );
  DFFRX1 \block_w2_reg_reg[2]  ( .D(n1325), .CK(clk), .RN(n1375), .Q(
        new_block[34]), .QN(n80) );
  DFFRX1 \block_w2_reg_reg[3]  ( .D(n1324), .CK(clk), .RN(n1376), .Q(
        new_block[35]), .QN(n79) );
  DFFRX1 \block_w3_reg_reg[0]  ( .D(n1359), .CK(clk), .RN(n1374), .Q(
        new_block[0]), .QN(n44) );
  DFFRX1 \block_w3_reg_reg[2]  ( .D(n1357), .CK(clk), .RN(n1375), .Q(
        new_block[2]), .QN(n42) );
  DFFRX1 \block_w3_reg_reg[3]  ( .D(n1356), .CK(clk), .RN(n1376), .Q(
        new_block[3]), .QN(n41) );
  DFFRX1 \block_w0_reg_reg[0]  ( .D(n1360), .CK(clk), .RN(n1373), .Q(
        new_block[96]), .QN(n146) );
  DFFRX1 \block_w0_reg_reg[14]  ( .D(n1250), .CK(clk), .RN(n1380), .Q(
        new_block[110]), .QN(n132) );
  DFFRX1 \block_w3_reg_reg[14]  ( .D(n1345), .CK(clk), .RN(n1379), .Q(
        new_block[14]), .QN(n30) );
  DFFRX1 \block_w1_reg_reg[12]  ( .D(n1283), .CK(clk), .RN(n1379), .Q(
        new_block[76]), .QN(n102) );
  DFFRX1 \block_w2_reg_reg[12]  ( .D(n1315), .CK(clk), .RN(n1376), .Q(
        new_block[44]), .QN(n70) );
  DFFRX1 \block_w1_reg_reg[10]  ( .D(n1285), .CK(clk), .RN(n1379), .Q(
        new_block[74]), .QN(n104) );
  DFFRX1 \block_w1_reg_reg[13]  ( .D(n1282), .CK(clk), .RN(n1379), .Q(
        new_block[77]), .QN(n101) );
  DFFRX1 \block_w1_reg_reg[14]  ( .D(n1281), .CK(clk), .RN(n1379), .Q(
        new_block[78]), .QN(n100) );
  DFFRX1 \block_w2_reg_reg[14]  ( .D(n1313), .CK(clk), .RN(n1380), .Q(
        new_block[46]), .QN(n68) );
  DFFRX1 \block_w2_reg_reg[13]  ( .D(n1314), .CK(clk), .RN(n1371), .Q(
        new_block[45]), .QN(n69) );
  DFFRX1 \block_w0_reg_reg[13]  ( .D(n1251), .CK(clk), .RN(n1372), .Q(
        new_block[109]), .QN(n133) );
  DFFRX1 \block_w3_reg_reg[13]  ( .D(n1346), .CK(clk), .RN(n1379), .Q(
        new_block[13]), .QN(n31) );
  DFFRX1 \block_w1_reg_reg[8]  ( .D(n1287), .CK(clk), .RN(n1378), .Q(
        new_block[72]), .QN(n106) );
  DFFRX1 \block_w1_reg_reg[9]  ( .D(n1286), .CK(clk), .RN(n1378), .Q(
        new_block[73]), .QN(n105) );
  DFFRX1 \block_w1_reg_reg[11]  ( .D(n1284), .CK(clk), .RN(n1379), .Q(
        new_block[75]), .QN(n103) );
  DFFRX1 \block_w2_reg_reg[9]  ( .D(n1318), .CK(clk), .RN(n1374), .Q(
        new_block[41]), .QN(n73) );
  DFFRX1 \block_w3_reg_reg[8]  ( .D(n1351), .CK(clk), .RN(n1378), .Q(
        new_block[8]), .QN(n36) );
  DFFRX1 \block_w3_reg_reg[9]  ( .D(n1350), .CK(clk), .RN(n1378), .Q(
        new_block[9]), .QN(n35) );
  DFFRX1 \block_w2_reg_reg[10]  ( .D(n1317), .CK(clk), .RN(n1375), .Q(
        new_block[42]), .QN(n72) );
  DFFRX1 \block_w0_reg_reg[10]  ( .D(n1254), .CK(clk), .RN(n1375), .Q(
        new_block[106]), .QN(n136) );
  DFFRX1 \block_w3_reg_reg[10]  ( .D(n1349), .CK(clk), .RN(n1378), .Q(
        new_block[10]), .QN(n34) );
  DFFRX1 \block_w2_reg_reg[8]  ( .D(n1319), .CK(clk), .RN(n1374), .Q(
        new_block[40]), .QN(n74) );
  DFFRX1 \block_w2_reg_reg[11]  ( .D(n1316), .CK(clk), .RN(n1375), .Q(
        new_block[43]), .QN(n71) );
  DFFRX1 \block_w3_reg_reg[12]  ( .D(n1347), .CK(clk), .RN(n1379), .Q(
        new_block[12]), .QN(n32) );
  DFFRX1 \block_w0_reg_reg[8]  ( .D(n1256), .CK(clk), .RN(n1374), .Q(
        new_block[104]), .QN(n138) );
  DFFRX1 \block_w0_reg_reg[12]  ( .D(n1252), .CK(clk), .RN(n1376), .Q(
        new_block[108]), .QN(n134) );
  DFFRX1 \block_w0_reg_reg[9]  ( .D(n1255), .CK(clk), .RN(n1374), .Q(
        new_block[105]), .QN(n137) );
  DFFRX1 \block_w0_reg_reg[11]  ( .D(n1253), .CK(clk), .RN(n1375), .Q(
        new_block[107]), .QN(n135) );
  DFFRX1 \block_w3_reg_reg[11]  ( .D(n1348), .CK(clk), .RN(n1379), .Q(
        new_block[11]), .QN(n33) );
  DFFRX1 \sword_ctr_reg_reg[1]  ( .D(n1368), .CK(clk), .RN(n1373), .Q(
        sword_ctr_reg[1]), .QN(n49) );
  DFFRX1 \sword_ctr_reg_reg[0]  ( .D(n1369), .CK(clk), .RN(n1373), .Q(
        sword_ctr_reg[0]), .QN(n50) );
  DFFRX1 \enc_ctrl_reg_reg[0]  ( .D(n1366), .CK(clk), .RN(n1373), .Q(
        enc_ctrl_reg[0]), .QN(n12) );
  DFFRX1 \round_ctr_reg_reg[3]  ( .D(n1362), .CK(clk), .RN(n1373), .Q(round[3]), .QN(n45) );
  DFFRX1 \round_ctr_reg_reg[2]  ( .D(n1363), .CK(clk), .RN(n1373), .Q(round[2]), .QN(n46) );
  DFFRX1 \enc_ctrl_reg_reg[1]  ( .D(n1367), .CK(clk), .RN(n1373), .Q(
        enc_ctrl_reg[1]), .QN(n11) );
  DFFRX1 \round_ctr_reg_reg[1]  ( .D(n1364), .CK(clk), .RN(n1373), .Q(round[1]), .QN(n47) );
  OAI221XL U3 ( .A0(n1224), .A1(n35), .B0(n218), .B1(n137), .C0(n221), .Y(
        sboxw[9]) );
  OA22X1 U4 ( .A0(n213), .A1(n104), .B0(n210), .B1(n72), .Y(n253) );
  OAI221XL U5 ( .A0(n256), .A1(n33), .B0(n218), .B1(n135), .C0(n252), .Y(
        sboxw[11]) );
  OA22X1 U6 ( .A0(n213), .A1(n103), .B0(n210), .B1(n71), .Y(n252) );
  OAI221XL U7 ( .A0(n256), .A1(n32), .B0(n218), .B1(n134), .C0(n251), .Y(
        sboxw[12]) );
  OA22X1 U8 ( .A0(n213), .A1(n102), .B0(n210), .B1(n70), .Y(n251) );
  NAND2X1 U9 ( .A(n969), .B(n728), .Y(n223) );
  OAI221XL U10 ( .A0(n1224), .A1(n36), .B0(n218), .B1(n138), .C0(n224), .Y(
        sboxw[8]) );
  OA22X1 U11 ( .A0(n215), .A1(n106), .B0(n212), .B1(n74), .Y(n224) );
  OA21XL U12 ( .A0(n1217), .A1(n1218), .B0(n1219), .Y(n1216) );
  OAI22XL U13 ( .A0(enc_ctrl_reg[1]), .A1(n1431), .B0(n1217), .B1(n1218), .Y(
        n1215) );
  NOR2X1 U14 ( .A(n1215), .B(n1216), .Y(n728) );
  NOR2X1 U15 ( .A(n1429), .B(n1216), .Y(n258) );
  OA21XL U16 ( .A0(keylen), .A1(n47), .B0(n46), .Y(n1229) );
  AOI211XL U17 ( .A0(n47), .A1(keylen), .B0(n1229), .C0(n45), .Y(n1217) );
  NAND2XL U18 ( .A(n12), .B(enc_ctrl_reg[1]), .Y(n1219) );
  NAND2X1 U19 ( .A(n730), .B(n728), .Y(n222) );
  NAND3XL U20 ( .A(n50), .B(n49), .C(n728), .Y(n220) );
  NAND2XL U21 ( .A(n729), .B(n256), .Y(n971) );
  NAND2XL U22 ( .A(n729), .B(n213), .Y(n491) );
  NAND2XL U23 ( .A(n729), .B(n220), .Y(n1) );
  NAND2XL U24 ( .A(n1431), .B(n1219), .Y(n1230) );
  NAND2XL U25 ( .A(n1431), .B(n1220), .Y(n1227) );
  OA22XL U26 ( .A0(n213), .A1(n101), .B0(n210), .B1(n69), .Y(n250) );
  OA22XL U27 ( .A0(n215), .A1(n105), .B0(n212), .B1(n73), .Y(n221) );
  OA22XL U28 ( .A0(n213), .A1(n100), .B0(n210), .B1(n68), .Y(n249) );
  OA22XL U29 ( .A0(n213), .A1(n114), .B0(n210), .B1(n82), .Y(n254) );
  OA22XL U30 ( .A0(n213), .A1(n99), .B0(n210), .B1(n67), .Y(n248) );
  OAI211XL U31 ( .A0(n1208), .A1(n1219), .B0(n1232), .C0(n1431), .Y(
        enc_ctrl_we) );
  NOR2XL U32 ( .A(n48), .B(n1431), .Y(n1223) );
  OAI21XL U33 ( .A0(n45), .A1(n2), .B0(n1222), .Y(n1362) );
  OA21XL U34 ( .A0(round[2]), .A1(n1431), .B0(n1225), .Y(n2) );
  NAND2BXL U35 ( .AN(n1208), .B(n728), .Y(n219) );
  NAND2XL U36 ( .A(n728), .B(n207), .Y(n255) );
  NAND2XL U37 ( .A(n728), .B(n155), .Y(n490) );
  BUFX2 U38 ( .A(n1381), .Y(n1380) );
  BUFX2 U39 ( .A(n1381), .Y(n1379) );
  BUFX2 U40 ( .A(n1382), .Y(n1378) );
  BUFX2 U41 ( .A(n1382), .Y(n1377) );
  BUFX2 U42 ( .A(n1383), .Y(n1376) );
  BUFX2 U43 ( .A(n1383), .Y(n1375) );
  BUFX2 U44 ( .A(n1384), .Y(n1374) );
  BUFX2 U45 ( .A(n1384), .Y(n1373) );
  BUFX2 U46 ( .A(n1371), .Y(n1381) );
  BUFX2 U47 ( .A(n1371), .Y(n1382) );
  BUFX2 U48 ( .A(n1371), .Y(n1383) );
  BUFX2 U49 ( .A(reset_n), .Y(n1370) );
  BUFX2 U50 ( .A(reset_n), .Y(n1371) );
  BUFX2 U51 ( .A(n1372), .Y(n1384) );
  BUFX2 U52 ( .A(reset_n), .Y(n1372) );
  NOR3BXL U53 ( .AN(n262), .B(n258), .C(n328), .Y(n729) );
  BUFX2 U54 ( .A(n732), .Y(n152) );
  BUFX2 U55 ( .A(n491), .Y(n155) );
  BUFX2 U56 ( .A(n1426), .Y(n7) );
  BUFX2 U57 ( .A(n1425), .Y(n6) );
  BUFX2 U58 ( .A(n1428), .Y(n148) );
  BUFX2 U59 ( .A(n209), .Y(n207) );
  BUFX2 U60 ( .A(n1425), .Y(n5) );
  BUFX2 U61 ( .A(n1428), .Y(n147) );
  BUFX2 U62 ( .A(n1426), .Y(n8) );
  INVX1 U63 ( .A(n166), .Y(n158) );
  INVX1 U64 ( .A(n166), .Y(n160) );
  INVX1 U65 ( .A(n166), .Y(n159) );
  INVX1 U66 ( .A(n165), .Y(n161) );
  INVX1 U67 ( .A(n175), .Y(n163) );
  INVX1 U68 ( .A(n165), .Y(n162) );
  BUFX2 U69 ( .A(n732), .Y(n154) );
  BUFX2 U70 ( .A(n732), .Y(n153) );
  BUFX2 U71 ( .A(n491), .Y(n157) );
  BUFX2 U72 ( .A(n491), .Y(n156) );
  BUFX2 U73 ( .A(n971), .Y(n149) );
  BUFX2 U74 ( .A(n1427), .Y(n10) );
  BUFX2 U75 ( .A(n971), .Y(n151) );
  BUFX2 U76 ( .A(n971), .Y(n150) );
  BUFX2 U77 ( .A(n1427), .Y(n9) );
  BUFX2 U78 ( .A(n209), .Y(n208) );
  BUFX2 U79 ( .A(n205), .Y(n193) );
  BUFX2 U80 ( .A(n203), .Y(n199) );
  BUFX2 U81 ( .A(n204), .Y(n196) );
  BUFX2 U82 ( .A(n205), .Y(n194) );
  BUFX2 U83 ( .A(n202), .Y(n200) );
  BUFX2 U84 ( .A(n203), .Y(n198) );
  BUFX2 U85 ( .A(n204), .Y(n197) );
  BUFX2 U86 ( .A(n202), .Y(n195) );
  BUFX2 U87 ( .A(n202), .Y(n201) );
  INVX1 U88 ( .A(n255), .Y(n1426) );
  INVX1 U89 ( .A(n731), .Y(n1428) );
  INVX1 U90 ( .A(n490), .Y(n1425) );
  BUFX2 U91 ( .A(n1), .Y(n209) );
  BUFX2 U92 ( .A(n175), .Y(n165) );
  BUFX2 U93 ( .A(n175), .Y(n166) );
  INVX1 U94 ( .A(n970), .Y(n1427) );
  BUFX2 U95 ( .A(n192), .Y(n176) );
  BUFX2 U96 ( .A(n192), .Y(n177) );
  INVX1 U97 ( .A(n165), .Y(n164) );
  BUFX2 U98 ( .A(n258), .Y(n206) );
  BUFX2 U99 ( .A(n258), .Y(n205) );
  BUFX2 U100 ( .A(n258), .Y(n202) );
  BUFX2 U101 ( .A(n258), .Y(n203) );
  BUFX2 U102 ( .A(n258), .Y(n204) );
  BUFX2 U103 ( .A(n173), .Y(n172) );
  BUFX2 U104 ( .A(n174), .Y(n167) );
  BUFX2 U105 ( .A(n173), .Y(n170) );
  BUFX2 U106 ( .A(n174), .Y(n169) );
  BUFX2 U107 ( .A(n174), .Y(n168) );
  BUFX2 U108 ( .A(n173), .Y(n171) );
  BUFX2 U109 ( .A(n188), .Y(n185) );
  BUFX2 U110 ( .A(n190), .Y(n181) );
  BUFX2 U111 ( .A(n191), .Y(n178) );
  BUFX2 U112 ( .A(n188), .Y(n184) );
  BUFX2 U113 ( .A(n189), .Y(n182) );
  BUFX2 U114 ( .A(n190), .Y(n180) );
  BUFX2 U115 ( .A(n189), .Y(n183) );
  BUFX2 U116 ( .A(n187), .Y(n186) );
  BUFX2 U117 ( .A(n191), .Y(n179) );
  BUFX2 U118 ( .A(n219), .Y(n256) );
  BUFX2 U119 ( .A(n223), .Y(n210) );
  BUFX2 U120 ( .A(n223), .Y(n212) );
  BUFX2 U121 ( .A(n222), .Y(n213) );
  BUFX2 U122 ( .A(n219), .Y(n1224) );
  BUFX2 U123 ( .A(n222), .Y(n215) );
  BUFX2 U124 ( .A(n223), .Y(n211) );
  BUFX2 U125 ( .A(n219), .Y(n1221) );
  BUFX2 U126 ( .A(n222), .Y(n214) );
  INVX1 U127 ( .A(new_sboxw[28]), .Y(n1388) );
  INVX1 U128 ( .A(new_sboxw[30]), .Y(n1395) );
  INVX1 U129 ( .A(new_sboxw[25]), .Y(n1389) );
  INVX1 U130 ( .A(new_sboxw[24]), .Y(n1390) );
  INVX1 U131 ( .A(new_sboxw[29]), .Y(n1393) );
  INVX1 U132 ( .A(new_sboxw[27]), .Y(n1392) );
  INVX1 U133 ( .A(new_sboxw[31]), .Y(n1394) );
  NAND2X1 U134 ( .A(n728), .B(n152), .Y(n731) );
  INVX1 U135 ( .A(new_sboxw[26]), .Y(n1391) );
  NAND2X1 U136 ( .A(n728), .B(n149), .Y(n970) );
  BUFX2 U137 ( .A(n262), .Y(n192) );
  BUFX2 U138 ( .A(n328), .Y(n175) );
  BUFX2 U139 ( .A(n328), .Y(n173) );
  BUFX2 U140 ( .A(n328), .Y(n174) );
  BUFX2 U141 ( .A(n262), .Y(n190) );
  BUFX2 U142 ( .A(n262), .Y(n188) );
  BUFX2 U143 ( .A(n262), .Y(n189) );
  BUFX2 U144 ( .A(n262), .Y(n191) );
  BUFX2 U145 ( .A(n262), .Y(n187) );
  BUFX2 U146 ( .A(n220), .Y(n218) );
  BUFX2 U147 ( .A(n220), .Y(n217) );
  BUFX2 U148 ( .A(n220), .Y(n216) );
  INVX1 U149 ( .A(n1215), .Y(n1429) );
  XOR2X1 U150 ( .A(n978), .B(n979), .Y(n977) );
  XOR2X1 U151 ( .A(n265), .B(n266), .Y(n264) );
  XOR2X1 U152 ( .A(n498), .B(n499), .Y(n497) );
  XOR2X1 U153 ( .A(n739), .B(n740), .Y(n738) );
  XOR2X1 U154 ( .A(n506), .B(n507), .Y(n505) );
  XOR2X1 U155 ( .A(n514), .B(n515), .Y(n513) );
  XOR2X1 U156 ( .A(n764), .B(n799), .Y(n798) );
  XOR2X1 U157 ( .A(n1003), .B(n1038), .Y(n1037) );
  XOR2X1 U158 ( .A(n273), .B(n274), .Y(n272) );
  XOR2X1 U159 ( .A(n281), .B(n282), .Y(n280) );
  XOR2X1 U160 ( .A(n308), .B(n309), .Y(n307) );
  XOR2X1 U161 ( .A(n747), .B(n748), .Y(n746) );
  XOR2X1 U162 ( .A(n755), .B(n756), .Y(n754) );
  XOR2X1 U163 ( .A(n782), .B(n783), .Y(n781) );
  XOR2X1 U164 ( .A(n986), .B(n987), .Y(n985) );
  XOR2X1 U165 ( .A(n290), .B(n325), .Y(n324) );
  XOR2X1 U166 ( .A(n523), .B(n558), .Y(n557) );
  XOR2X1 U167 ( .A(n994), .B(n995), .Y(n993) );
  XOR2X1 U168 ( .A(n1021), .B(n1022), .Y(n1020) );
  XOR2X1 U169 ( .A(n541), .B(n542), .Y(n540) );
  NAND2BX1 U170 ( .AN(n1219), .B(enc_ctrl_we), .Y(n1228) );
  INVX1 U171 ( .A(n1223), .Y(n1430) );
  NOR2X1 U172 ( .A(n50), .B(sword_ctr_reg[1]), .Y(n730) );
  NOR2X1 U173 ( .A(n49), .B(sword_ctr_reg[0]), .Y(n969) );
  OAI221XL U174 ( .A0(n256), .A1(n34), .B0(n218), .B1(n136), .C0(n253), .Y(
        sboxw[10]) );
  OAI221XL U175 ( .A0(n256), .A1(n30), .B0(n218), .B1(n132), .C0(n249), .Y(
        sboxw[14]) );
  INVX1 U176 ( .A(enc_ctrl_reg[0]), .Y(n1431) );
  OAI221XL U177 ( .A0(n256), .A1(n31), .B0(n218), .B1(n133), .C0(n250), .Y(
        sboxw[13]) );
  NAND2X1 U178 ( .A(enc_ctrl_reg[0]), .B(enc_ctrl_reg[1]), .Y(n1218) );
  NAND2X1 U179 ( .A(sword_ctr_reg[1]), .B(sword_ctr_reg[0]), .Y(n1208) );
  OAI221XL U180 ( .A0(n256), .A1(n29), .B0(n218), .B1(n131), .C0(n248), .Y(
        sboxw[15]) );
  OAI221XL U181 ( .A0(n256), .A1(n44), .B0(n218), .B1(n146), .C0(n254), .Y(
        sboxw[0]) );
  OAI221XL U182 ( .A0(n1221), .A1(n42), .B0(n217), .B1(n144), .C0(n232), .Y(
        sboxw[2]) );
  OA22X1 U183 ( .A0(n215), .A1(n112), .B0(n211), .B1(n80), .Y(n232) );
  OAI221XL U184 ( .A0(n1221), .A1(n39), .B0(n217), .B1(n141), .C0(n227), .Y(
        sboxw[5]) );
  OA22X1 U185 ( .A0(n215), .A1(n109), .B0(n211), .B1(n77), .Y(n227) );
  OA22X1 U186 ( .A0(n215), .A1(n110), .B0(n211), .B1(n78), .Y(n228) );
  NAND3X1 U187 ( .A(n3), .B(n4), .C(n228), .Y(sboxw[4]) );
  OR2X1 U188 ( .A(n217), .B(n142), .Y(n4) );
  OAI221XL U189 ( .A0(n1224), .A1(n43), .B0(n216), .B1(n145), .C0(n243), .Y(
        sboxw[1]) );
  OAI221XL U190 ( .A0(n1221), .A1(n41), .B0(n217), .B1(n143), .C0(n229), .Y(
        sboxw[3]) );
  OA22X1 U191 ( .A0(n215), .A1(n111), .B0(n211), .B1(n79), .Y(n229) );
  OA22X1 U192 ( .A0(n214), .A1(n113), .B0(n212), .B1(n81), .Y(n243) );
  OAI221XL U193 ( .A0(n644), .A1(n180), .B0(n103), .B1(n156), .C0(n645), .Y(
        n1284) );
  XNOR2X1 U194 ( .A(round_key[75]), .B(block[75]), .Y(n644) );
  AOI222XL U195 ( .A0(n6), .A1(new_sboxw[11]), .B0(n169), .B1(n646), .C0(n197), 
        .C1(n647), .Y(n645) );
  XOR2X1 U196 ( .A(round_key[75]), .B(new_block[11]), .Y(n646) );
  OAI221XL U197 ( .A0(n1124), .A1(n185), .B0(n33), .B1(n150), .C0(n1125), .Y(
        n1348) );
  XNOR2X1 U198 ( .A(round_key[11]), .B(block[11]), .Y(n1124) );
  AOI222XL U199 ( .A0(n10), .A1(new_sboxw[11]), .B0(n174), .B1(n1126), .C0(
        n195), .C1(n1127), .Y(n1125) );
  XOR2X1 U200 ( .A(round_key[11]), .B(new_block[75]), .Y(n1126) );
  OAI221XL U201 ( .A0(n885), .A1(n178), .B0(n71), .B1(n153), .C0(n886), .Y(
        n1316) );
  XNOR2X1 U202 ( .A(round_key[43]), .B(block[43]), .Y(n885) );
  AOI222XL U203 ( .A0(n148), .A1(new_sboxw[11]), .B0(n167), .B1(n887), .C0(
        n200), .C1(n888), .Y(n886) );
  XOR2X1 U204 ( .A(round_key[43]), .B(new_block[107]), .Y(n887) );
  OAI221XL U205 ( .A0(n412), .A1(n184), .B0(n135), .B1(n208), .C0(n413), .Y(
        n1253) );
  XNOR2X1 U206 ( .A(round_key[107]), .B(block[107]), .Y(n412) );
  AOI222XL U207 ( .A0(new_sboxw[11]), .A1(n7), .B0(n171), .B1(n414), .C0(n203), 
        .C1(n415), .Y(n413) );
  XOR2X1 U208 ( .A(round_key[107]), .B(new_block[43]), .Y(n414) );
  OAI221XL U209 ( .A0(n1221), .A1(n38), .B0(n217), .B1(n140), .C0(n226), .Y(
        sboxw[6]) );
  OA22X1 U210 ( .A0(n222), .A1(n108), .B0(n211), .B1(n76), .Y(n226) );
  OAI221XL U211 ( .A0(n1224), .A1(n37), .B0(n218), .B1(n139), .C0(n225), .Y(
        sboxw[7]) );
  OAI221XL U212 ( .A0(n445), .A1(n183), .B0(n140), .B1(n207), .C0(n446), .Y(
        n1258) );
  XNOR2X1 U213 ( .A(round_key[102]), .B(block[102]), .Y(n445) );
  XOR2X1 U214 ( .A(round_key[102]), .B(new_block[6]), .Y(n447) );
  OAI221XL U215 ( .A0(n1202), .A1(n186), .B0(n44), .B1(n149), .C0(n1203), .Y(
        n1359) );
  XNOR2X1 U216 ( .A(round_key[0]), .B(block[0]), .Y(n1202) );
  AOI222XL U217 ( .A0(n9), .A1(new_sboxw[0]), .B0(n165), .B1(n1204), .C0(n193), 
        .C1(n1205), .Y(n1203) );
  XOR2X1 U218 ( .A(round_key[0]), .B(new_block[32]), .Y(n1204) );
  OAI221XL U219 ( .A0(n963), .A1(n182), .B0(n82), .B1(n152), .C0(n964), .Y(
        n1327) );
  XNOR2X1 U220 ( .A(round_key[32]), .B(block[32]), .Y(n963) );
  AOI222XL U221 ( .A0(n147), .A1(new_sboxw[0]), .B0(n166), .B1(n965), .C0(n201), .C1(n966), .Y(n964) );
  XOR2X1 U222 ( .A(round_key[32]), .B(new_block[64]), .Y(n965) );
  OAI221XL U223 ( .A0(n722), .A1(n179), .B0(n114), .B1(n155), .C0(n723), .Y(
        n1295) );
  XNOR2X1 U224 ( .A(round_key[64]), .B(block[64]), .Y(n722) );
  AOI222XL U225 ( .A0(new_sboxw[0]), .A1(n5), .B0(n168), .B1(n724), .C0(n198), 
        .C1(n725), .Y(n723) );
  XOR2X1 U226 ( .A(round_key[64]), .B(new_block[96]), .Y(n724) );
  OAI221XL U227 ( .A0(n1209), .A1(n187), .B0(n146), .B1(n207), .C0(n1210), .Y(
        n1360) );
  XNOR2X1 U228 ( .A(round_key[96]), .B(block[96]), .Y(n1209) );
  AOI222XL U229 ( .A0(new_sboxw[0]), .A1(n1426), .B0(n175), .B1(n1211), .C0(
        n197), .C1(n1212), .Y(n1210) );
  OAI221XL U230 ( .A0(n1221), .A1(n15), .B0(n217), .B1(n117), .C0(n233), .Y(
        sboxw[29]) );
  OAI221XL U231 ( .A0(n1221), .A1(n16), .B0(n217), .B1(n118), .C0(n234), .Y(
        sboxw[28]) );
  OAI221XL U232 ( .A0(n1221), .A1(n17), .B0(n217), .B1(n119), .C0(n235), .Y(
        sboxw[27]) );
  OAI221XL U233 ( .A0(n1224), .A1(n20), .B0(n216), .B1(n122), .C0(n238), .Y(
        sboxw[24]) );
  OAI221XL U234 ( .A0(n1224), .A1(n19), .B0(n216), .B1(n121), .C0(n237), .Y(
        sboxw[25]) );
  OAI221XL U235 ( .A0(n871), .A1(n178), .B0(n69), .B1(n153), .C0(n872), .Y(
        n1314) );
  XNOR2X1 U236 ( .A(round_key[45]), .B(block[45]), .Y(n871) );
  AOI222XL U237 ( .A0(n148), .A1(new_sboxw[13]), .B0(n167), .B1(n873), .C0(
        n200), .C1(n874), .Y(n872) );
  XOR2X1 U238 ( .A(round_key[45]), .B(new_block[109]), .Y(n873) );
  OAI221XL U239 ( .A0(n630), .A1(n180), .B0(n101), .B1(n156), .C0(n631), .Y(
        n1282) );
  XNOR2X1 U240 ( .A(round_key[77]), .B(block[77]), .Y(n630) );
  AOI222XL U241 ( .A0(n6), .A1(new_sboxw[13]), .B0(n169), .B1(n632), .C0(n197), 
        .C1(n633), .Y(n631) );
  XOR2X1 U242 ( .A(round_key[77]), .B(new_block[13]), .Y(n632) );
  OAI221XL U243 ( .A0(n1110), .A1(n185), .B0(n31), .B1(n150), .C0(n1111), .Y(
        n1346) );
  XNOR2X1 U244 ( .A(round_key[13]), .B(block[13]), .Y(n1110) );
  AOI222XL U245 ( .A0(n10), .A1(new_sboxw[13]), .B0(n174), .B1(n1112), .C0(
        n196), .C1(n1113), .Y(n1111) );
  XOR2X1 U246 ( .A(round_key[13]), .B(new_block[77]), .Y(n1112) );
  OAI221XL U247 ( .A0(n1157), .A1(n186), .B0(n38), .B1(n149), .C0(n1158), .Y(
        n1353) );
  XNOR2X1 U248 ( .A(round_key[6]), .B(block[6]), .Y(n1157) );
  XOR2X1 U249 ( .A(round_key[6]), .B(new_block[38]), .Y(n1159) );
  OAI221XL U250 ( .A0(n918), .A1(n181), .B0(n76), .B1(n152), .C0(n919), .Y(
        n1321) );
  XNOR2X1 U251 ( .A(round_key[38]), .B(block[38]), .Y(n918) );
  XOR2X1 U252 ( .A(round_key[38]), .B(new_block[70]), .Y(n920) );
  OAI221XL U253 ( .A0(n677), .A1(n179), .B0(n108), .B1(n155), .C0(n678), .Y(
        n1289) );
  XNOR2X1 U254 ( .A(round_key[70]), .B(block[70]), .Y(n677) );
  XOR2X1 U255 ( .A(round_key[70]), .B(new_block[102]), .Y(n679) );
  OAI221XL U256 ( .A0(n256), .A1(n28), .B0(n220), .B1(n130), .C0(n247), .Y(
        sboxw[16]) );
  OAI221XL U257 ( .A0(n256), .A1(n27), .B0(n220), .B1(n129), .C0(n246), .Y(
        sboxw[17]) );
  OAI221XL U258 ( .A0(n859), .A1(n178), .B0(n67), .B1(n153), .C0(n860), .Y(
        n1312) );
  XNOR2X1 U259 ( .A(round_key[47]), .B(block[47]), .Y(n859) );
  AOI222XL U260 ( .A0(n148), .A1(new_sboxw[15]), .B0(n167), .B1(n861), .C0(
        n200), .C1(n862), .Y(n860) );
  XOR2X1 U261 ( .A(round_key[47]), .B(new_block[111]), .Y(n861) );
  OAI221XL U262 ( .A0(n670), .A1(n179), .B0(n107), .B1(n155), .C0(n671), .Y(
        n1288) );
  XNOR2X1 U263 ( .A(round_key[71]), .B(block[71]), .Y(n670) );
  AOI222XL U264 ( .A0(n5), .A1(new_sboxw[7]), .B0(n169), .B1(n672), .C0(n197), 
        .C1(n673), .Y(n671) );
  XOR2X1 U265 ( .A(round_key[71]), .B(new_block[103]), .Y(n672) );
  OAI221XL U266 ( .A0(n1098), .A1(n183), .B0(n29), .B1(n150), .C0(n1099), .Y(
        n1344) );
  XNOR2X1 U267 ( .A(round_key[15]), .B(block[15]), .Y(n1098) );
  AOI222XL U268 ( .A0(n10), .A1(new_sboxw[15]), .B0(n166), .B1(n1100), .C0(
        n198), .C1(n1101), .Y(n1099) );
  XOR2X1 U269 ( .A(round_key[15]), .B(new_block[79]), .Y(n1100) );
  OAI221XL U270 ( .A0(n911), .A1(n179), .B0(n75), .B1(n152), .C0(n912), .Y(
        n1320) );
  XNOR2X1 U271 ( .A(round_key[39]), .B(block[39]), .Y(n911) );
  AOI222XL U272 ( .A0(n147), .A1(new_sboxw[7]), .B0(n174), .B1(n913), .C0(n201), .C1(n914), .Y(n912) );
  XOR2X1 U273 ( .A(round_key[39]), .B(new_block[71]), .Y(n913) );
  OAI221XL U274 ( .A0(n1150), .A1(n186), .B0(n37), .B1(n149), .C0(n1151), .Y(
        n1352) );
  XNOR2X1 U275 ( .A(round_key[7]), .B(block[7]), .Y(n1150) );
  AOI222XL U276 ( .A0(n9), .A1(new_sboxw[7]), .B0(n173), .B1(n1152), .C0(n195), 
        .C1(n1153), .Y(n1151) );
  XOR2X1 U277 ( .A(round_key[7]), .B(new_block[39]), .Y(n1152) );
  OAI221XL U278 ( .A0(n618), .A1(n180), .B0(n99), .B1(n156), .C0(n619), .Y(
        n1280) );
  XNOR2X1 U279 ( .A(round_key[79]), .B(block[79]), .Y(n618) );
  AOI222XL U280 ( .A0(n6), .A1(new_sboxw[15]), .B0(n169), .B1(n620), .C0(n197), 
        .C1(n621), .Y(n619) );
  XOR2X1 U281 ( .A(round_key[79]), .B(new_block[15]), .Y(n620) );
  OAI221XL U282 ( .A0(n438), .A1(n183), .B0(n139), .B1(n207), .C0(n439), .Y(
        n1257) );
  XNOR2X1 U283 ( .A(round_key[103]), .B(block[103]), .Y(n438) );
  AOI222XL U284 ( .A0(new_sboxw[7]), .A1(n8), .B0(n171), .B1(n440), .C0(n203), 
        .C1(n441), .Y(n439) );
  XOR2X1 U285 ( .A(round_key[103]), .B(new_block[7]), .Y(n440) );
  XNOR2X1 U286 ( .A(round_key[76]), .B(block[76]), .Y(n636) );
  XOR2X1 U287 ( .A(round_key[76]), .B(new_block[12]), .Y(n638) );
  XNOR2X1 U288 ( .A(round_key[12]), .B(block[12]), .Y(n1116) );
  XOR2X1 U289 ( .A(round_key[12]), .B(new_block[76]), .Y(n1118) );
  XNOR2X1 U290 ( .A(round_key[44]), .B(block[44]), .Y(n877) );
  XOR2X1 U291 ( .A(round_key[44]), .B(new_block[108]), .Y(n879) );
  XNOR2X1 U292 ( .A(round_key[72]), .B(block[72]), .Y(n664) );
  XOR2X1 U293 ( .A(round_key[72]), .B(new_block[8]), .Y(n666) );
  XNOR2X1 U294 ( .A(round_key[8]), .B(block[8]), .Y(n1144) );
  XOR2X1 U295 ( .A(round_key[8]), .B(new_block[72]), .Y(n1146) );
  XNOR2X1 U296 ( .A(round_key[4]), .B(block[4]), .Y(n1171) );
  XOR2X1 U297 ( .A(round_key[4]), .B(new_block[36]), .Y(n1173) );
  XNOR2X1 U298 ( .A(round_key[36]), .B(block[36]), .Y(n932) );
  XOR2X1 U299 ( .A(round_key[36]), .B(new_block[68]), .Y(n934) );
  XNOR2X1 U300 ( .A(round_key[68]), .B(block[68]), .Y(n691) );
  XOR2X1 U301 ( .A(round_key[68]), .B(new_block[100]), .Y(n693) );
  XNOR2X1 U302 ( .A(round_key[100]), .B(block[100]), .Y(n459) );
  XOR2X1 U303 ( .A(round_key[100]), .B(new_block[4]), .Y(n461) );
  XNOR2X1 U304 ( .A(round_key[108]), .B(block[108]), .Y(n404) );
  XOR2X1 U305 ( .A(round_key[108]), .B(new_block[44]), .Y(n406) );
  XNOR2X1 U306 ( .A(round_key[1]), .B(block[1]), .Y(n1194) );
  XOR2X1 U307 ( .A(round_key[1]), .B(new_block[33]), .Y(n1196) );
  XNOR2X1 U308 ( .A(round_key[33]), .B(block[33]), .Y(n955) );
  XOR2X1 U309 ( .A(round_key[33]), .B(new_block[65]), .Y(n957) );
  XNOR2X1 U310 ( .A(round_key[65]), .B(block[65]), .Y(n714) );
  XOR2X1 U311 ( .A(round_key[65]), .B(new_block[97]), .Y(n716) );
  XNOR2X1 U312 ( .A(round_key[97]), .B(block[97]), .Y(n482) );
  XOR2X1 U313 ( .A(round_key[97]), .B(new_block[1]), .Y(n484) );
  XNOR2X1 U314 ( .A(round_key[40]), .B(block[40]), .Y(n905) );
  XOR2X1 U315 ( .A(round_key[40]), .B(new_block[104]), .Y(n907) );
  XNOR2X1 U316 ( .A(round_key[104]), .B(block[104]), .Y(n432) );
  XOR2X1 U317 ( .A(round_key[104]), .B(new_block[40]), .Y(n434) );
  OAI221XL U318 ( .A0(n1221), .A1(n14), .B0(n217), .B1(n116), .C0(n231), .Y(
        sboxw[30]) );
  OAI221XL U319 ( .A0(n1395), .A1(n731), .B0(n52), .B1(n732), .C0(n741), .Y(
        n1297) );
  AOI222XL U320 ( .A0(n202), .A1(n742), .B0(n743), .B1(n1411), .C0(
        round_key[62]), .C1(n744), .Y(n741) );
  INVX1 U321 ( .A(round_key[62]), .Y(n1411) );
  XOR2X1 U322 ( .A(n745), .B(n746), .Y(n742) );
  OAI221XL U323 ( .A0(n1054), .A1(n182), .B0(n23), .B1(n151), .C0(n1055), .Y(
        n1338) );
  XNOR2X1 U324 ( .A(round_key[21]), .B(block[21]), .Y(n1054) );
  AOI222XL U325 ( .A0(n1427), .A1(new_sboxw[21]), .B0(n173), .B1(n1056), .C0(
        n199), .C1(n1057), .Y(n1055) );
  XOR2X1 U326 ( .A(round_key[21]), .B(new_block[117]), .Y(n1056) );
  OAI221XL U327 ( .A0(n1393), .A1(n970), .B0(n15), .B1(n971), .C0(n988), .Y(
        n1330) );
  AOI222XL U328 ( .A0(n202), .A1(n989), .B0(n990), .B1(n1416), .C0(
        round_key[29]), .C1(n991), .Y(n988) );
  INVX1 U329 ( .A(round_key[29]), .Y(n1416) );
  XOR2X1 U330 ( .A(n992), .B(n993), .Y(n989) );
  OAI221XL U331 ( .A0(n349), .A1(n185), .B0(n126), .B1(n209), .C0(n350), .Y(
        n1244) );
  XNOR2X1 U332 ( .A(round_key[116]), .B(block[116]), .Y(n349) );
  AOI222XL U333 ( .A0(new_sboxw[20]), .A1(n8), .B0(n172), .B1(n351), .C0(n194), 
        .C1(n352), .Y(n350) );
  XOR2X1 U334 ( .A(round_key[116]), .B(new_block[84]), .Y(n351) );
  OAI221XL U335 ( .A0(n581), .A1(n181), .B0(n94), .B1(n157), .C0(n582), .Y(
        n1275) );
  XNOR2X1 U336 ( .A(round_key[84]), .B(block[84]), .Y(n581) );
  AOI222XL U337 ( .A0(n1425), .A1(new_sboxw[20]), .B0(n170), .B1(n583), .C0(
        n196), .C1(n584), .Y(n582) );
  XOR2X1 U338 ( .A(round_key[84]), .B(new_block[52]), .Y(n583) );
  OAI221XL U339 ( .A0(n822), .A1(n189), .B0(n62), .B1(n154), .C0(n823), .Y(
        n1307) );
  XNOR2X1 U340 ( .A(round_key[52]), .B(block[52]), .Y(n822) );
  AOI222XL U341 ( .A0(n1428), .A1(new_sboxw[20]), .B0(n167), .B1(n824), .C0(
        n199), .C1(n825), .Y(n823) );
  XOR2X1 U342 ( .A(round_key[52]), .B(new_block[20]), .Y(n824) );
  OAI221XL U343 ( .A0(n1061), .A1(n182), .B0(n24), .B1(n151), .C0(n1062), .Y(
        n1339) );
  XNOR2X1 U344 ( .A(round_key[20]), .B(block[20]), .Y(n1061) );
  AOI222XL U345 ( .A0(n1427), .A1(new_sboxw[20]), .B0(n165), .B1(n1063), .C0(
        n199), .C1(n1064), .Y(n1062) );
  XOR2X1 U346 ( .A(round_key[20]), .B(new_block[116]), .Y(n1063) );
  OAI221XL U347 ( .A0(n1388), .A1(n970), .B0(n16), .B1(n151), .C0(n996), .Y(
        n1331) );
  AOI222XL U348 ( .A0(n202), .A1(n997), .B0(n998), .B1(n1420), .C0(
        round_key[28]), .C1(n999), .Y(n996) );
  INVX1 U349 ( .A(round_key[28]), .Y(n1420) );
  OAI22XL U350 ( .A0(n16), .A1(n158), .B0(n192), .B1(n1451), .Y(n998) );
  OAI221XL U351 ( .A0(n357), .A1(n185), .B0(n127), .B1(n209), .C0(n358), .Y(
        n1245) );
  XNOR2X1 U352 ( .A(round_key[115]), .B(block[115]), .Y(n357) );
  AOI222XL U353 ( .A0(new_sboxw[19]), .A1(n7), .B0(n172), .B1(n359), .C0(n194), 
        .C1(n360), .Y(n358) );
  XOR2X1 U354 ( .A(round_key[115]), .B(new_block[83]), .Y(n359) );
  OAI221XL U355 ( .A0(n589), .A1(n181), .B0(n95), .B1(n157), .C0(n590), .Y(
        n1276) );
  XNOR2X1 U356 ( .A(round_key[83]), .B(block[83]), .Y(n589) );
  AOI222XL U357 ( .A0(n6), .A1(new_sboxw[19]), .B0(n170), .B1(n591), .C0(n196), 
        .C1(n592), .Y(n590) );
  XOR2X1 U358 ( .A(round_key[83]), .B(new_block[51]), .Y(n591) );
  OAI221XL U359 ( .A0(n830), .A1(n187), .B0(n63), .B1(n154), .C0(n831), .Y(
        n1308) );
  XNOR2X1 U360 ( .A(round_key[51]), .B(block[51]), .Y(n830) );
  AOI222XL U361 ( .A0(n148), .A1(new_sboxw[19]), .B0(n167), .B1(n832), .C0(
        n199), .C1(n833), .Y(n831) );
  XOR2X1 U362 ( .A(round_key[51]), .B(new_block[19]), .Y(n832) );
  OAI221XL U363 ( .A0(n1069), .A1(n182), .B0(n25), .B1(n151), .C0(n1070), .Y(
        n1340) );
  XNOR2X1 U364 ( .A(round_key[19]), .B(block[19]), .Y(n1069) );
  AOI222XL U365 ( .A0(n10), .A1(new_sboxw[19]), .B0(n166), .B1(n1071), .C0(
        n199), .C1(n1072), .Y(n1070) );
  XOR2X1 U366 ( .A(round_key[19]), .B(new_block[115]), .Y(n1071) );
  OAI221XL U367 ( .A0(n1392), .A1(n970), .B0(n17), .B1(n151), .C0(n1006), .Y(
        n1332) );
  AOI222XL U368 ( .A0(n203), .A1(n1007), .B0(n1008), .B1(n1408), .C0(
        round_key[27]), .C1(n1009), .Y(n1006) );
  INVX1 U369 ( .A(round_key[27]), .Y(n1408) );
  OAI22XL U370 ( .A0(n17), .A1(n158), .B0(n192), .B1(n1447), .Y(n1008) );
  OAI221XL U371 ( .A0(n365), .A1(n184), .B0(n128), .B1(n208), .C0(n366), .Y(
        n1246) );
  XNOR2X1 U372 ( .A(round_key[114]), .B(block[114]), .Y(n365) );
  AOI222XL U373 ( .A0(new_sboxw[18]), .A1(n7), .B0(n172), .B1(n367), .C0(n194), 
        .C1(n368), .Y(n366) );
  XOR2X1 U374 ( .A(round_key[114]), .B(new_block[82]), .Y(n367) );
  OAI221XL U375 ( .A0(n597), .A1(n181), .B0(n96), .B1(n156), .C0(n598), .Y(
        n1277) );
  XNOR2X1 U376 ( .A(round_key[82]), .B(block[82]), .Y(n597) );
  AOI222XL U377 ( .A0(n6), .A1(new_sboxw[18]), .B0(n170), .B1(n599), .C0(n196), 
        .C1(n600), .Y(n598) );
  XOR2X1 U378 ( .A(round_key[82]), .B(new_block[50]), .Y(n599) );
  OAI221XL U379 ( .A0(n838), .A1(n178), .B0(n64), .B1(n153), .C0(n839), .Y(
        n1309) );
  XNOR2X1 U380 ( .A(round_key[50]), .B(block[50]), .Y(n838) );
  AOI222XL U381 ( .A0(n148), .A1(new_sboxw[18]), .B0(n167), .B1(n840), .C0(
        n200), .C1(n841), .Y(n839) );
  XOR2X1 U382 ( .A(round_key[50]), .B(new_block[18]), .Y(n840) );
  OAI221XL U383 ( .A0(n1077), .A1(n182), .B0(n26), .B1(n150), .C0(n1078), .Y(
        n1341) );
  XNOR2X1 U384 ( .A(round_key[18]), .B(block[18]), .Y(n1077) );
  AOI222XL U385 ( .A0(n10), .A1(new_sboxw[18]), .B0(n166), .B1(n1079), .C0(
        n199), .C1(n1080), .Y(n1078) );
  XOR2X1 U386 ( .A(round_key[18]), .B(new_block[114]), .Y(n1079) );
  OAI221XL U387 ( .A0(n604), .A1(n180), .B0(n97), .B1(n156), .C0(n605), .Y(
        n1278) );
  XNOR2X1 U388 ( .A(round_key[81]), .B(block[81]), .Y(n604) );
  AOI222XL U389 ( .A0(n6), .A1(new_sboxw[17]), .B0(n170), .B1(n606), .C0(n196), 
        .C1(n607), .Y(n605) );
  XOR2X1 U390 ( .A(round_key[81]), .B(new_block[49]), .Y(n606) );
  OAI221XL U391 ( .A0(n845), .A1(n178), .B0(n65), .B1(n153), .C0(n846), .Y(
        n1310) );
  XNOR2X1 U392 ( .A(round_key[49]), .B(block[49]), .Y(n845) );
  AOI222XL U393 ( .A0(n148), .A1(new_sboxw[17]), .B0(n167), .B1(n847), .C0(
        n200), .C1(n848), .Y(n846) );
  XOR2X1 U394 ( .A(round_key[49]), .B(new_block[17]), .Y(n847) );
  OAI221XL U395 ( .A0(n1084), .A1(n182), .B0(n27), .B1(n150), .C0(n1085), .Y(
        n1342) );
  XNOR2X1 U396 ( .A(round_key[17]), .B(block[17]), .Y(n1084) );
  AOI222XL U397 ( .A0(n10), .A1(new_sboxw[17]), .B0(n165), .B1(n1086), .C0(
        n198), .C1(n1087), .Y(n1085) );
  XOR2X1 U398 ( .A(round_key[17]), .B(new_block[113]), .Y(n1086) );
  OAI221XL U399 ( .A0(n1389), .A1(n970), .B0(n19), .B1(n151), .C0(n1023), .Y(
        n1334) );
  AOI222XL U400 ( .A0(n193), .A1(n1024), .B0(n1025), .B1(n1424), .C0(
        round_key[25]), .C1(n1026), .Y(n1023) );
  INVX1 U401 ( .A(round_key[25]), .Y(n1424) );
  OAI22XL U402 ( .A0(n19), .A1(n158), .B0(n176), .B1(n1434), .Y(n1025) );
  OAI221XL U403 ( .A0(n372), .A1(n184), .B0(n129), .B1(n208), .C0(n373), .Y(
        n1247) );
  XNOR2X1 U404 ( .A(round_key[113]), .B(block[113]), .Y(n372) );
  AOI222XL U405 ( .A0(new_sboxw[17]), .A1(n7), .B0(n172), .B1(n374), .C0(n194), 
        .C1(n375), .Y(n373) );
  XOR2X1 U406 ( .A(round_key[113]), .B(new_block[81]), .Y(n374) );
  OAI221XL U407 ( .A0(n612), .A1(n180), .B0(n98), .B1(n156), .C0(n613), .Y(
        n1279) );
  XNOR2X1 U408 ( .A(round_key[80]), .B(block[80]), .Y(n612) );
  AOI222XL U409 ( .A0(n6), .A1(new_sboxw[16]), .B0(n169), .B1(n614), .C0(n196), 
        .C1(n615), .Y(n613) );
  XOR2X1 U410 ( .A(round_key[80]), .B(new_block[48]), .Y(n614) );
  OAI221XL U411 ( .A0(n853), .A1(n178), .B0(n66), .B1(n153), .C0(n854), .Y(
        n1311) );
  XNOR2X1 U412 ( .A(round_key[48]), .B(block[48]), .Y(n853) );
  AOI222XL U413 ( .A0(n148), .A1(new_sboxw[16]), .B0(n167), .B1(n855), .C0(
        n200), .C1(n856), .Y(n854) );
  XOR2X1 U414 ( .A(round_key[48]), .B(new_block[16]), .Y(n855) );
  OAI221XL U415 ( .A0(n1390), .A1(n731), .B0(n58), .B1(n154), .C0(n793), .Y(
        n1303) );
  AOI222XL U416 ( .A0(n204), .A1(n794), .B0(n795), .B1(n1399), .C0(
        round_key[56]), .C1(n796), .Y(n793) );
  INVX1 U417 ( .A(round_key[56]), .Y(n1399) );
  XOR2X1 U418 ( .A(n797), .B(n798), .Y(n794) );
  OAI221XL U419 ( .A0(n335), .A1(n185), .B0(n124), .B1(n209), .C0(n336), .Y(
        n1242) );
  XNOR2X1 U420 ( .A(round_key[118]), .B(block[118]), .Y(n335) );
  AOI222XL U421 ( .A0(new_sboxw[22]), .A1(n8), .B0(n172), .B1(n337), .C0(n194), 
        .C1(n338), .Y(n336) );
  XOR2X1 U422 ( .A(round_key[118]), .B(new_block[86]), .Y(n337) );
  OAI221XL U423 ( .A0(n574), .A1(n181), .B0(n93), .B1(n157), .C0(n575), .Y(
        n1274) );
  XNOR2X1 U424 ( .A(round_key[85]), .B(block[85]), .Y(n574) );
  AOI222XL U425 ( .A0(n1425), .A1(new_sboxw[21]), .B0(n170), .B1(n576), .C0(
        n196), .C1(n577), .Y(n575) );
  XOR2X1 U426 ( .A(round_key[85]), .B(new_block[53]), .Y(n576) );
  OAI221XL U427 ( .A0(n815), .A1(n191), .B0(n61), .B1(n154), .C0(n816), .Y(
        n1306) );
  XNOR2X1 U428 ( .A(round_key[53]), .B(block[53]), .Y(n815) );
  AOI222XL U429 ( .A0(n1428), .A1(new_sboxw[21]), .B0(n168), .B1(n817), .C0(
        n199), .C1(n818), .Y(n816) );
  XOR2X1 U430 ( .A(round_key[53]), .B(new_block[21]), .Y(n817) );
  OAI221XL U431 ( .A0(n1393), .A1(n731), .B0(n53), .B1(n732), .C0(n749), .Y(
        n1298) );
  AOI222XL U432 ( .A0(n204), .A1(n750), .B0(n751), .B1(n1415), .C0(
        round_key[61]), .C1(n752), .Y(n749) );
  INVX1 U433 ( .A(round_key[61]), .Y(n1415) );
  XOR2X1 U434 ( .A(n753), .B(n754), .Y(n750) );
  OAI221XL U435 ( .A0(n1388), .A1(n731), .B0(n54), .B1(n154), .C0(n757), .Y(
        n1299) );
  AOI222XL U436 ( .A0(n205), .A1(n758), .B0(n759), .B1(n1419), .C0(
        round_key[60]), .C1(n760), .Y(n757) );
  INVX1 U437 ( .A(round_key[60]), .Y(n1419) );
  OAI22XL U438 ( .A0(n54), .A1(n160), .B0(n192), .B1(n1450), .Y(n759) );
  OAI221XL U439 ( .A0(n1392), .A1(n731), .B0(n55), .B1(n154), .C0(n767), .Y(
        n1300) );
  AOI222XL U440 ( .A0(n205), .A1(n768), .B0(n769), .B1(n1407), .C0(
        round_key[59]), .C1(n770), .Y(n767) );
  INVX1 U441 ( .A(round_key[59]), .Y(n1407) );
  OAI22XL U442 ( .A0(n55), .A1(n159), .B0(n192), .B1(n1446), .Y(n769) );
  OAI221XL U443 ( .A0(n1389), .A1(n731), .B0(n57), .B1(n154), .C0(n784), .Y(
        n1302) );
  AOI222XL U444 ( .A0(n202), .A1(n785), .B0(n786), .B1(n1423), .C0(
        round_key[57]), .C1(n787), .Y(n784) );
  INVX1 U445 ( .A(round_key[57]), .Y(n1423) );
  OAI22XL U446 ( .A0(n57), .A1(n159), .B0(n188), .B1(n1432), .Y(n786) );
  OAI221XL U447 ( .A0(n1092), .A1(n183), .B0(n28), .B1(n150), .C0(n1093), .Y(
        n1343) );
  XNOR2X1 U448 ( .A(round_key[16]), .B(block[16]), .Y(n1092) );
  AOI222XL U449 ( .A0(n10), .A1(new_sboxw[16]), .B0(n165), .B1(n1094), .C0(
        n198), .C1(n1095), .Y(n1093) );
  XOR2X1 U450 ( .A(round_key[16]), .B(new_block[112]), .Y(n1094) );
  OAI221XL U451 ( .A0(n1390), .A1(n970), .B0(n20), .B1(n151), .C0(n1032), .Y(
        n1335) );
  AOI222XL U452 ( .A0(n193), .A1(n1033), .B0(n1034), .B1(n1400), .C0(
        round_key[24]), .C1(n1035), .Y(n1032) );
  INVX1 U453 ( .A(round_key[24]), .Y(n1400) );
  XOR2X1 U454 ( .A(n1036), .B(n1037), .Y(n1033) );
  OAI221XL U455 ( .A0(n1394), .A1(n970), .B0(n13), .B1(n971), .C0(n972), .Y(
        n1328) );
  AOI222XL U456 ( .A0(n203), .A1(n973), .B0(n974), .B1(n1396), .C0(
        round_key[31]), .C1(n975), .Y(n972) );
  INVX1 U457 ( .A(round_key[31]), .Y(n1396) );
  XOR2X1 U458 ( .A(n976), .B(n977), .Y(n973) );
  OAI221XL U459 ( .A0(n1395), .A1(n970), .B0(n14), .B1(n971), .C0(n980), .Y(
        n1329) );
  AOI222XL U460 ( .A0(n204), .A1(n981), .B0(n982), .B1(n1412), .C0(
        round_key[30]), .C1(n983), .Y(n980) );
  INVX1 U461 ( .A(round_key[30]), .Y(n1412) );
  XOR2X1 U462 ( .A(n984), .B(n985), .Y(n981) );
  OAI221XL U463 ( .A0(n342), .A1(n185), .B0(n125), .B1(n209), .C0(n343), .Y(
        n1243) );
  XNOR2X1 U464 ( .A(round_key[117]), .B(block[117]), .Y(n342) );
  AOI222XL U465 ( .A0(new_sboxw[21]), .A1(n8), .B0(n172), .B1(n344), .C0(n194), 
        .C1(n345), .Y(n343) );
  XOR2X1 U466 ( .A(round_key[117]), .B(new_block[85]), .Y(n344) );
  OAI221XL U467 ( .A0(n398), .A1(n184), .B0(n133), .B1(n208), .C0(n399), .Y(
        n1251) );
  XNOR2X1 U468 ( .A(round_key[109]), .B(block[109]), .Y(n398) );
  AOI222XL U469 ( .A0(new_sboxw[13]), .A1(n7), .B0(n171), .B1(n400), .C0(n202), 
        .C1(n401), .Y(n399) );
  XOR2X1 U470 ( .A(round_key[109]), .B(new_block[45]), .Y(n400) );
  OAI221XL U471 ( .A0(n255), .A1(n1395), .B0(n116), .B1(n208), .C0(n267), .Y(
        n1234) );
  AOI222XL U472 ( .A0(n206), .A1(n268), .B0(n269), .B1(n1409), .C0(
        round_key[126]), .C1(n270), .Y(n267) );
  INVX1 U473 ( .A(round_key[126]), .Y(n1409) );
  XOR2X1 U474 ( .A(n271), .B(n272), .Y(n268) );
  OAI221XL U475 ( .A0(n255), .A1(n1393), .B0(n117), .B1(n208), .C0(n275), .Y(
        n1235) );
  AOI222XL U476 ( .A0(n206), .A1(n276), .B0(n277), .B1(n1413), .C0(
        round_key[125]), .C1(n278), .Y(n275) );
  INVX1 U477 ( .A(round_key[125]), .Y(n1413) );
  XOR2X1 U478 ( .A(n279), .B(n280), .Y(n276) );
  OAI221XL U479 ( .A0(n255), .A1(n1388), .B0(n118), .B1(n1), .C0(n283), .Y(
        n1236) );
  AOI222XL U480 ( .A0(n206), .A1(n284), .B0(n285), .B1(n1417), .C0(
        round_key[124]), .C1(n286), .Y(n283) );
  INVX1 U481 ( .A(round_key[124]), .Y(n1417) );
  OAI22XL U482 ( .A0(n118), .A1(n159), .B0(n189), .B1(n1448), .Y(n285) );
  OAI221XL U483 ( .A0(n255), .A1(n1392), .B0(n119), .B1(n1), .C0(n293), .Y(
        n1237) );
  AOI222XL U484 ( .A0(n206), .A1(n294), .B0(n295), .B1(n1405), .C0(
        round_key[123]), .C1(n296), .Y(n293) );
  INVX1 U485 ( .A(round_key[123]), .Y(n1405) );
  OAI22XL U486 ( .A0(n119), .A1(n159), .B0(n191), .B1(n1444), .Y(n295) );
  OAI221XL U487 ( .A0(n255), .A1(n1389), .B0(n121), .B1(n1), .C0(n310), .Y(
        n1239) );
  AOI222XL U488 ( .A0(n206), .A1(n311), .B0(n312), .B1(n1421), .C0(
        round_key[121]), .C1(n313), .Y(n310) );
  INVX1 U489 ( .A(round_key[121]), .Y(n1421) );
  OAI22XL U490 ( .A0(n121), .A1(n160), .B0(n188), .B1(n1433), .Y(n312) );
  OAI221XL U491 ( .A0(n255), .A1(n1390), .B0(n122), .B1(n1), .C0(n319), .Y(
        n1240) );
  AOI222XL U492 ( .A0(n206), .A1(n320), .B0(n321), .B1(n1397), .C0(
        round_key[120]), .C1(n322), .Y(n319) );
  INVX1 U493 ( .A(round_key[120]), .Y(n1397) );
  XOR2X1 U494 ( .A(n323), .B(n324), .Y(n320) );
  OAI221XL U495 ( .A0(n255), .A1(n1394), .B0(n115), .B1(n208), .C0(n257), .Y(
        n1233) );
  AOI222XL U496 ( .A0(n202), .A1(n259), .B0(n260), .B1(n1385), .C0(
        round_key[127]), .C1(n261), .Y(n257) );
  INVX1 U497 ( .A(round_key[127]), .Y(n1385) );
  XOR2X1 U498 ( .A(n263), .B(n264), .Y(n259) );
  OAI221XL U499 ( .A0(n567), .A1(n181), .B0(n92), .B1(n157), .C0(n568), .Y(
        n1273) );
  XNOR2X1 U500 ( .A(round_key[86]), .B(block[86]), .Y(n567) );
  AOI222XL U501 ( .A0(n1425), .A1(new_sboxw[22]), .B0(n170), .B1(n569), .C0(
        n196), .C1(n570), .Y(n568) );
  XOR2X1 U502 ( .A(round_key[86]), .B(new_block[54]), .Y(n569) );
  OAI221XL U503 ( .A0(n1395), .A1(n490), .B0(n84), .B1(n491), .C0(n500), .Y(
        n1265) );
  AOI222XL U504 ( .A0(n206), .A1(n501), .B0(n502), .B1(n1410), .C0(
        round_key[94]), .C1(n503), .Y(n500) );
  INVX1 U505 ( .A(round_key[94]), .Y(n1410) );
  XOR2X1 U506 ( .A(n504), .B(n505), .Y(n501) );
  OAI221XL U507 ( .A0(n1393), .A1(n490), .B0(n85), .B1(n491), .C0(n508), .Y(
        n1266) );
  AOI222XL U508 ( .A0(n203), .A1(n509), .B0(n510), .B1(n1414), .C0(
        round_key[93]), .C1(n511), .Y(n508) );
  INVX1 U509 ( .A(round_key[93]), .Y(n1414) );
  XOR2X1 U510 ( .A(n512), .B(n513), .Y(n509) );
  OAI221XL U511 ( .A0(n1388), .A1(n490), .B0(n86), .B1(n157), .C0(n516), .Y(
        n1267) );
  AOI222XL U512 ( .A0(n204), .A1(n517), .B0(n518), .B1(n1418), .C0(
        round_key[92]), .C1(n519), .Y(n516) );
  INVX1 U513 ( .A(round_key[92]), .Y(n1418) );
  OAI22XL U514 ( .A0(n86), .A1(n160), .B0(n187), .B1(n1449), .Y(n518) );
  OAI221XL U515 ( .A0(n1392), .A1(n490), .B0(n87), .B1(n157), .C0(n526), .Y(
        n1268) );
  AOI222XL U516 ( .A0(n205), .A1(n527), .B0(n528), .B1(n1406), .C0(
        round_key[91]), .C1(n529), .Y(n526) );
  INVX1 U517 ( .A(round_key[91]), .Y(n1406) );
  OAI22XL U518 ( .A0(n87), .A1(n161), .B0(n176), .B1(n1445), .Y(n528) );
  OAI221XL U519 ( .A0(n1389), .A1(n490), .B0(n89), .B1(n157), .C0(n543), .Y(
        n1270) );
  AOI222XL U520 ( .A0(n204), .A1(n544), .B0(n545), .B1(n1422), .C0(
        round_key[89]), .C1(n546), .Y(n543) );
  INVX1 U521 ( .A(round_key[89]), .Y(n1422) );
  OAI22XL U522 ( .A0(n89), .A1(n160), .B0(n187), .B1(n1435), .Y(n545) );
  OAI221XL U523 ( .A0(n1390), .A1(n490), .B0(n90), .B1(n157), .C0(n552), .Y(
        n1271) );
  AOI222XL U524 ( .A0(n205), .A1(n553), .B0(n554), .B1(n1398), .C0(
        round_key[88]), .C1(n555), .Y(n552) );
  INVX1 U525 ( .A(round_key[88]), .Y(n1398) );
  XOR2X1 U526 ( .A(n556), .B(n557), .Y(n553) );
  OAI221XL U527 ( .A0(n1394), .A1(n490), .B0(n83), .B1(n491), .C0(n492), .Y(
        n1264) );
  AOI222XL U528 ( .A0(n206), .A1(n493), .B0(n494), .B1(n1386), .C0(
        round_key[95]), .C1(n495), .Y(n492) );
  INVX1 U529 ( .A(round_key[95]), .Y(n1386) );
  XOR2X1 U530 ( .A(n496), .B(n497), .Y(n493) );
  OAI221XL U531 ( .A0(n808), .A1(n190), .B0(n60), .B1(n154), .C0(n809), .Y(
        n1305) );
  XNOR2X1 U532 ( .A(round_key[54]), .B(block[54]), .Y(n808) );
  AOI222XL U533 ( .A0(n1428), .A1(new_sboxw[22]), .B0(n168), .B1(n810), .C0(
        n199), .C1(n811), .Y(n809) );
  XOR2X1 U534 ( .A(round_key[54]), .B(new_block[22]), .Y(n810) );
  OAI221XL U535 ( .A0(n392), .A1(n184), .B0(n132), .B1(n208), .C0(n393), .Y(
        n1250) );
  XNOR2X1 U536 ( .A(round_key[110]), .B(block[110]), .Y(n392) );
  AOI222XL U537 ( .A0(new_sboxw[14]), .A1(n7), .B0(n172), .B1(n394), .C0(n202), 
        .C1(n395), .Y(n393) );
  XOR2X1 U538 ( .A(round_key[110]), .B(new_block[46]), .Y(n394) );
  OAI221XL U539 ( .A0(n865), .A1(n178), .B0(n68), .B1(n153), .C0(n866), .Y(
        n1313) );
  XNOR2X1 U540 ( .A(round_key[46]), .B(block[46]), .Y(n865) );
  AOI222XL U541 ( .A0(n148), .A1(new_sboxw[14]), .B0(n167), .B1(n867), .C0(
        n200), .C1(n868), .Y(n866) );
  XOR2X1 U542 ( .A(round_key[46]), .B(new_block[110]), .Y(n867) );
  OAI221XL U543 ( .A0(n1394), .A1(n731), .B0(n51), .B1(n732), .C0(n733), .Y(
        n1296) );
  AOI222XL U544 ( .A0(n203), .A1(n734), .B0(n735), .B1(n1387), .C0(
        round_key[63]), .C1(n736), .Y(n733) );
  INVX1 U545 ( .A(round_key[63]), .Y(n1387) );
  XOR2X1 U546 ( .A(n737), .B(n738), .Y(n734) );
  OAI221XL U547 ( .A0(n1047), .A1(n182), .B0(n22), .B1(n151), .C0(n1048), .Y(
        n1337) );
  XNOR2X1 U548 ( .A(round_key[22]), .B(block[22]), .Y(n1047) );
  AOI222XL U549 ( .A0(n1427), .A1(new_sboxw[22]), .B0(n165), .B1(n1049), .C0(
        n199), .C1(n1050), .Y(n1048) );
  XOR2X1 U550 ( .A(round_key[22]), .B(new_block[118]), .Y(n1049) );
  OAI221XL U551 ( .A0(n624), .A1(n180), .B0(n100), .B1(n156), .C0(n625), .Y(
        n1281) );
  XNOR2X1 U552 ( .A(round_key[78]), .B(block[78]), .Y(n624) );
  AOI222XL U553 ( .A0(n6), .A1(new_sboxw[14]), .B0(n169), .B1(n626), .C0(n197), 
        .C1(n627), .Y(n625) );
  XOR2X1 U554 ( .A(round_key[78]), .B(new_block[14]), .Y(n626) );
  OAI221XL U555 ( .A0(n1104), .A1(n185), .B0(n30), .B1(n150), .C0(n1105), .Y(
        n1345) );
  XNOR2X1 U556 ( .A(round_key[14]), .B(block[14]), .Y(n1104) );
  AOI222XL U557 ( .A0(n10), .A1(new_sboxw[14]), .B0(n174), .B1(n1106), .C0(
        n196), .C1(n1107), .Y(n1105) );
  XOR2X1 U558 ( .A(round_key[14]), .B(new_block[78]), .Y(n1106) );
  OAI221XL U559 ( .A0(n651), .A1(n180), .B0(n104), .B1(n156), .C0(n652), .Y(
        n1285) );
  XNOR2X1 U560 ( .A(round_key[74]), .B(block[74]), .Y(n651) );
  AOI222XL U561 ( .A0(n6), .A1(new_sboxw[10]), .B0(n169), .B1(n653), .C0(n197), 
        .C1(n654), .Y(n652) );
  XOR2X1 U562 ( .A(round_key[74]), .B(new_block[10]), .Y(n653) );
  OAI221XL U563 ( .A0(n1131), .A1(n185), .B0(n34), .B1(n150), .C0(n1132), .Y(
        n1349) );
  XNOR2X1 U564 ( .A(round_key[10]), .B(block[10]), .Y(n1131) );
  AOI222XL U565 ( .A0(n10), .A1(new_sboxw[10]), .B0(n173), .B1(n1133), .C0(
        n195), .C1(n1134), .Y(n1132) );
  XOR2X1 U566 ( .A(round_key[10]), .B(new_block[74]), .Y(n1133) );
  OAI221XL U567 ( .A0(n657), .A1(n180), .B0(n105), .B1(n156), .C0(n658), .Y(
        n1286) );
  XNOR2X1 U568 ( .A(round_key[73]), .B(block[73]), .Y(n657) );
  XOR2X1 U569 ( .A(round_key[73]), .B(new_block[9]), .Y(n659) );
  OAI221XL U570 ( .A0(n1137), .A1(n186), .B0(n35), .B1(n150), .C0(n1138), .Y(
        n1350) );
  XNOR2X1 U571 ( .A(round_key[9]), .B(block[9]), .Y(n1137) );
  XOR2X1 U572 ( .A(round_key[9]), .B(new_block[73]), .Y(n1139) );
  OAI221XL U573 ( .A0(n380), .A1(n184), .B0(n130), .B1(n209), .C0(n381), .Y(
        n1248) );
  XNOR2X1 U574 ( .A(round_key[112]), .B(block[112]), .Y(n380) );
  AOI222XL U575 ( .A0(new_sboxw[16]), .A1(n7), .B0(n172), .B1(n382), .C0(n194), 
        .C1(n383), .Y(n381) );
  XOR2X1 U576 ( .A(round_key[112]), .B(new_block[80]), .Y(n382) );
  OAI221XL U577 ( .A0(n1164), .A1(n186), .B0(n39), .B1(n149), .C0(n1165), .Y(
        n1354) );
  XNOR2X1 U578 ( .A(round_key[5]), .B(block[5]), .Y(n1164) );
  AOI222XL U579 ( .A0(n9), .A1(new_sboxw[5]), .B0(n175), .B1(n1166), .C0(n193), 
        .C1(n1167), .Y(n1165) );
  XOR2X1 U580 ( .A(round_key[5]), .B(new_block[37]), .Y(n1166) );
  OAI221XL U581 ( .A0(n925), .A1(n181), .B0(n77), .B1(n152), .C0(n926), .Y(
        n1322) );
  XNOR2X1 U582 ( .A(round_key[37]), .B(block[37]), .Y(n925) );
  AOI222XL U583 ( .A0(n147), .A1(new_sboxw[5]), .B0(n173), .B1(n927), .C0(n201), .C1(n928), .Y(n926) );
  XOR2X1 U584 ( .A(round_key[37]), .B(new_block[69]), .Y(n927) );
  OAI221XL U585 ( .A0(n684), .A1(n179), .B0(n109), .B1(n155), .C0(n685), .Y(
        n1290) );
  XNOR2X1 U586 ( .A(round_key[69]), .B(block[69]), .Y(n684) );
  AOI222XL U587 ( .A0(n5), .A1(new_sboxw[5]), .B0(n168), .B1(n686), .C0(n198), 
        .C1(n687), .Y(n685) );
  XOR2X1 U588 ( .A(round_key[69]), .B(new_block[101]), .Y(n686) );
  OAI221XL U589 ( .A0(n892), .A1(n178), .B0(n72), .B1(n153), .C0(n893), .Y(
        n1317) );
  XNOR2X1 U590 ( .A(round_key[42]), .B(block[42]), .Y(n892) );
  AOI222XL U591 ( .A0(n148), .A1(new_sboxw[10]), .B0(n173), .B1(n894), .C0(
        n200), .C1(n895), .Y(n893) );
  XOR2X1 U592 ( .A(round_key[42]), .B(new_block[106]), .Y(n894) );
  OAI221XL U593 ( .A0(n1187), .A1(n186), .B0(n42), .B1(n149), .C0(n1188), .Y(
        n1357) );
  XNOR2X1 U594 ( .A(round_key[2]), .B(block[2]), .Y(n1187) );
  AOI222XL U595 ( .A0(n9), .A1(new_sboxw[2]), .B0(n165), .B1(n1189), .C0(n193), 
        .C1(n1190), .Y(n1188) );
  XOR2X1 U596 ( .A(round_key[2]), .B(new_block[34]), .Y(n1189) );
  OAI221XL U597 ( .A0(n948), .A1(n182), .B0(n80), .B1(n152), .C0(n949), .Y(
        n1325) );
  XNOR2X1 U598 ( .A(round_key[34]), .B(block[34]), .Y(n948) );
  AOI222XL U599 ( .A0(n147), .A1(new_sboxw[2]), .B0(n166), .B1(n950), .C0(n201), .C1(n951), .Y(n949) );
  XOR2X1 U600 ( .A(round_key[34]), .B(new_block[66]), .Y(n950) );
  OAI221XL U601 ( .A0(n707), .A1(n179), .B0(n112), .B1(n155), .C0(n708), .Y(
        n1293) );
  XNOR2X1 U602 ( .A(round_key[66]), .B(block[66]), .Y(n707) );
  AOI222XL U603 ( .A0(n5), .A1(new_sboxw[2]), .B0(n168), .B1(n709), .C0(n198), 
        .C1(n710), .Y(n708) );
  XOR2X1 U604 ( .A(round_key[66]), .B(new_block[98]), .Y(n709) );
  OAI221XL U605 ( .A0(n475), .A1(n183), .B0(n144), .B1(n207), .C0(n476), .Y(
        n1262) );
  XNOR2X1 U606 ( .A(round_key[98]), .B(block[98]), .Y(n475) );
  AOI222XL U607 ( .A0(new_sboxw[2]), .A1(n8), .B0(n170), .B1(n477), .C0(n195), 
        .C1(n478), .Y(n476) );
  XOR2X1 U608 ( .A(round_key[98]), .B(new_block[2]), .Y(n477) );
  OAI221XL U609 ( .A0(n898), .A1(n178), .B0(n73), .B1(n153), .C0(n899), .Y(
        n1318) );
  XNOR2X1 U610 ( .A(round_key[41]), .B(block[41]), .Y(n898) );
  XOR2X1 U611 ( .A(round_key[41]), .B(new_block[105]), .Y(n900) );
  OAI221XL U612 ( .A0(n425), .A1(n184), .B0(n137), .B1(n209), .C0(n426), .Y(
        n1255) );
  XNOR2X1 U613 ( .A(round_key[105]), .B(block[105]), .Y(n425) );
  XOR2X1 U614 ( .A(round_key[105]), .B(new_block[41]), .Y(n427) );
  OAI221XL U615 ( .A0(n1039), .A1(n182), .B0(n21), .B1(n151), .C0(n1040), .Y(
        n1336) );
  XNOR2X1 U616 ( .A(round_key[23]), .B(block[23]), .Y(n1039) );
  AOI222XL U617 ( .A0(n1427), .A1(new_sboxw[23]), .B0(n166), .B1(n1041), .C0(
        n193), .C1(n1042), .Y(n1040) );
  XOR2X1 U618 ( .A(round_key[23]), .B(new_block[119]), .Y(n1041) );
  OAI221XL U619 ( .A0(n386), .A1(n184), .B0(n131), .B1(n208), .C0(n387), .Y(
        n1249) );
  XNOR2X1 U620 ( .A(round_key[111]), .B(block[111]), .Y(n386) );
  AOI222XL U621 ( .A0(new_sboxw[15]), .A1(n7), .B0(n172), .B1(n388), .C0(n194), 
        .C1(n389), .Y(n387) );
  XOR2X1 U622 ( .A(round_key[111]), .B(new_block[47]), .Y(n388) );
  OAI221XL U623 ( .A0(n1179), .A1(n186), .B0(n41), .B1(n149), .C0(n1180), .Y(
        n1356) );
  XNOR2X1 U624 ( .A(round_key[3]), .B(block[3]), .Y(n1179) );
  AOI222XL U625 ( .A0(n9), .A1(new_sboxw[3]), .B0(n175), .B1(n1181), .C0(n193), 
        .C1(n1182), .Y(n1180) );
  XOR2X1 U626 ( .A(round_key[3]), .B(new_block[35]), .Y(n1181) );
  OAI221XL U627 ( .A0(n940), .A1(n181), .B0(n79), .B1(n152), .C0(n941), .Y(
        n1324) );
  XNOR2X1 U628 ( .A(round_key[35]), .B(block[35]), .Y(n940) );
  AOI222XL U629 ( .A0(n147), .A1(new_sboxw[3]), .B0(n175), .B1(n942), .C0(n201), .C1(n943), .Y(n941) );
  XOR2X1 U630 ( .A(round_key[35]), .B(new_block[67]), .Y(n942) );
  OAI221XL U631 ( .A0(n699), .A1(n179), .B0(n111), .B1(n155), .C0(n700), .Y(
        n1292) );
  XNOR2X1 U632 ( .A(round_key[67]), .B(block[67]), .Y(n699) );
  AOI222XL U633 ( .A0(n5), .A1(new_sboxw[3]), .B0(n168), .B1(n701), .C0(n198), 
        .C1(n702), .Y(n700) );
  XOR2X1 U634 ( .A(round_key[67]), .B(new_block[99]), .Y(n701) );
  OAI221XL U635 ( .A0(n467), .A1(n183), .B0(n143), .B1(n207), .C0(n468), .Y(
        n1261) );
  XNOR2X1 U636 ( .A(round_key[99]), .B(block[99]), .Y(n467) );
  AOI222XL U637 ( .A0(new_sboxw[3]), .A1(n1426), .B0(n170), .B1(n469), .C0(
        n195), .C1(n470), .Y(n468) );
  XOR2X1 U638 ( .A(round_key[99]), .B(new_block[3]), .Y(n469) );
  OAI221XL U639 ( .A0(n326), .A1(n185), .B0(n123), .B1(n209), .C0(n327), .Y(
        n1241) );
  XNOR2X1 U640 ( .A(round_key[119]), .B(block[119]), .Y(n326) );
  AOI222XL U641 ( .A0(new_sboxw[23]), .A1(n8), .B0(n172), .B1(n329), .C0(n194), 
        .C1(n330), .Y(n327) );
  XOR2X1 U642 ( .A(round_key[119]), .B(new_block[87]), .Y(n329) );
  OAI221XL U643 ( .A0(n559), .A1(n181), .B0(n91), .B1(n157), .C0(n560), .Y(
        n1272) );
  XNOR2X1 U644 ( .A(round_key[87]), .B(block[87]), .Y(n559) );
  AOI222XL U645 ( .A0(n1425), .A1(new_sboxw[23]), .B0(n170), .B1(n561), .C0(
        n196), .C1(n562), .Y(n560) );
  XOR2X1 U646 ( .A(round_key[87]), .B(new_block[55]), .Y(n561) );
  OAI221XL U647 ( .A0(n800), .A1(n188), .B0(n59), .B1(n154), .C0(n801), .Y(
        n1304) );
  XNOR2X1 U648 ( .A(round_key[55]), .B(block[55]), .Y(n800) );
  AOI222XL U649 ( .A0(n1428), .A1(new_sboxw[23]), .B0(n168), .B1(n802), .C0(
        n199), .C1(n803), .Y(n801) );
  XOR2X1 U650 ( .A(round_key[55]), .B(new_block[23]), .Y(n802) );
  OAI221XL U651 ( .A0(n452), .A1(n183), .B0(n141), .B1(n207), .C0(n453), .Y(
        n1259) );
  XNOR2X1 U652 ( .A(round_key[101]), .B(block[101]), .Y(n452) );
  AOI222XL U653 ( .A0(new_sboxw[5]), .A1(n1426), .B0(n171), .B1(n454), .C0(
        n204), .C1(n455), .Y(n453) );
  XOR2X1 U654 ( .A(round_key[101]), .B(new_block[5]), .Y(n454) );
  OAI221XL U655 ( .A0(n419), .A1(n184), .B0(n136), .B1(n209), .C0(n420), .Y(
        n1254) );
  XNOR2X1 U656 ( .A(round_key[106]), .B(block[106]), .Y(n419) );
  AOI222XL U657 ( .A0(new_sboxw[10]), .A1(n7), .B0(n171), .B1(n421), .C0(n205), 
        .C1(n422), .Y(n420) );
  XOR2X1 U658 ( .A(round_key[106]), .B(new_block[42]), .Y(n421) );
  OAI221XL U659 ( .A0(n1221), .A1(n13), .B0(n217), .B1(n115), .C0(n230), .Y(
        sboxw[31]) );
  OAI221XL U660 ( .A0(n1391), .A1(n970), .B0(n18), .B1(n151), .C0(n1015), .Y(
        n1333) );
  AOI222XL U661 ( .A0(n193), .A1(n1016), .B0(n1017), .B1(n1404), .C0(
        round_key[26]), .C1(n1018), .Y(n1015) );
  INVX1 U662 ( .A(round_key[26]), .Y(n1404) );
  XOR2X1 U663 ( .A(n1019), .B(n1020), .Y(n1016) );
  OAI221XL U664 ( .A0(n1391), .A1(n731), .B0(n56), .B1(n154), .C0(n776), .Y(
        n1301) );
  AOI222XL U665 ( .A0(n205), .A1(n777), .B0(n778), .B1(n1403), .C0(
        round_key[58]), .C1(n779), .Y(n776) );
  INVX1 U666 ( .A(round_key[58]), .Y(n1403) );
  XOR2X1 U667 ( .A(n780), .B(n781), .Y(n777) );
  OAI221XL U668 ( .A0(n255), .A1(n1391), .B0(n120), .B1(n208), .C0(n302), .Y(
        n1238) );
  AOI222XL U669 ( .A0(n206), .A1(n303), .B0(n304), .B1(n1401), .C0(
        round_key[122]), .C1(n305), .Y(n302) );
  INVX1 U670 ( .A(round_key[122]), .Y(n1401) );
  XOR2X1 U671 ( .A(n306), .B(n307), .Y(n303) );
  OAI221XL U672 ( .A0(n1391), .A1(n490), .B0(n88), .B1(n157), .C0(n535), .Y(
        n1269) );
  AOI222XL U673 ( .A0(n203), .A1(n536), .B0(n537), .B1(n1402), .C0(
        round_key[90]), .C1(n538), .Y(n535) );
  INVX1 U674 ( .A(round_key[90]), .Y(n1402) );
  XOR2X1 U675 ( .A(n539), .B(n540), .Y(n536) );
  XOR2X1 U676 ( .A(round_key[84]), .B(new_block[92]), .Y(n588) );
  XOR2X1 U677 ( .A(round_key[65]), .B(new_block[9]), .Y(n721) );
  XOR2X1 U678 ( .A(round_key[116]), .B(new_block[83]), .Y(n356) );
  XOR2X1 U679 ( .A(round_key[20]), .B(new_block[75]), .Y(n1068) );
  XOR2X1 U680 ( .A(round_key[115]), .B(new_block[82]), .Y(n364) );
  XOR2X1 U681 ( .A(round_key[19]), .B(new_block[74]), .Y(n1076) );
  XOR2X1 U682 ( .A(round_key[17]), .B(new_block[72]), .Y(n1091) );
  XOR2X1 U683 ( .A(round_key[113]), .B(new_block[80]), .Y(n379) );
  XOR2X1 U684 ( .A(round_key[4]), .B(new_block[76]), .Y(n1178) );
  XOR2X1 U685 ( .A(round_key[36]), .B(new_block[67]), .Y(n939) );
  XOR2X1 U686 ( .A(round_key[68]), .B(new_block[99]), .Y(n698) );
  XOR2X1 U687 ( .A(round_key[3]), .B(new_block[75]), .Y(n1186) );
  XOR2X1 U688 ( .A(round_key[35]), .B(new_block[66]), .Y(n947) );
  XOR2X1 U689 ( .A(round_key[67]), .B(new_block[98]), .Y(n706) );
  XOR2X1 U690 ( .A(round_key[1]), .B(new_block[73]), .Y(n1201) );
  XOR2X1 U691 ( .A(round_key[33]), .B(new_block[64]), .Y(n962) );
  XOR2X1 U692 ( .A(n1058), .B(n1059), .Y(n1057) );
  XOR2X1 U693 ( .A(new_block[116]), .B(n994), .Y(n1059) );
  XOR2X1 U694 ( .A(new_block[29]), .B(n1060), .Y(n1058) );
  XOR2X1 U695 ( .A(round_key[21]), .B(new_block[76]), .Y(n1060) );
  XOR2X1 U696 ( .A(n287), .B(n288), .Y(n284) );
  XOR2X1 U697 ( .A(n289), .B(n290), .Y(n288) );
  XOR2X1 U698 ( .A(n291), .B(n292), .Y(n287) );
  XOR2X1 U699 ( .A(round_key[124]), .B(new_block[84]), .Y(n292) );
  XOR2X1 U700 ( .A(n297), .B(n298), .Y(n294) );
  XOR2X1 U701 ( .A(n299), .B(n300), .Y(n298) );
  XOR2X1 U702 ( .A(n290), .B(n301), .Y(n297) );
  XOR2X1 U703 ( .A(round_key[123]), .B(new_block[83]), .Y(n301) );
  XOR2X1 U704 ( .A(n314), .B(n315), .Y(n311) );
  XOR2X1 U705 ( .A(n316), .B(n317), .Y(n315) );
  XOR2X1 U706 ( .A(n290), .B(n318), .Y(n314) );
  XOR2X1 U707 ( .A(round_key[121]), .B(new_block[81]), .Y(n318) );
  XOR2X1 U708 ( .A(n881), .B(n882), .Y(n880) );
  XOR2X1 U709 ( .A(n773), .B(n883), .Y(n882) );
  XOR2X1 U710 ( .A(n756), .B(n884), .Y(n881) );
  XOR2X1 U711 ( .A(round_key[44]), .B(new_block[68]), .Y(n884) );
  XOR2X1 U712 ( .A(n902), .B(n903), .Y(n901) );
  XOR2X1 U713 ( .A(n799), .B(n883), .Y(n903) );
  XOR2X1 U714 ( .A(n783), .B(n904), .Y(n902) );
  XOR2X1 U715 ( .A(round_key[41]), .B(new_block[65]), .Y(n904) );
  XOR2X1 U716 ( .A(round_key[52]), .B(new_block[60]), .Y(n829) );
  XOR2X1 U717 ( .A(round_key[49]), .B(new_block[57]), .Y(n852) );
  XOR2X1 U718 ( .A(round_key[81]), .B(new_block[8]), .Y(n611) );
  XOR2X1 U719 ( .A(round_key[97]), .B(new_block[41]), .Y(n489) );
  XOR2X1 U720 ( .A(round_key[100]), .B(new_block[44]), .Y(n466) );
  XOR2X1 U721 ( .A(round_key[83]), .B(new_block[91]), .Y(n596) );
  XOR2X1 U722 ( .A(round_key[51]), .B(new_block[59]), .Y(n837) );
  XOR2X1 U723 ( .A(round_key[99]), .B(new_block[43]), .Y(n474) );
  XOR2X1 U724 ( .A(n922), .B(n923), .Y(n921) );
  XOR2X1 U725 ( .A(new_block[110]), .B(n739), .Y(n923) );
  XOR2X1 U726 ( .A(new_block[61]), .B(n924), .Y(n922) );
  XOR2X1 U727 ( .A(round_key[38]), .B(new_block[69]), .Y(n924) );
  XOR2X1 U728 ( .A(n1175), .B(n1176), .Y(n1174) );
  XOR2X1 U729 ( .A(n1177), .B(n1045), .Y(n1176) );
  XOR2X1 U730 ( .A(n79), .B(n1178), .Y(n1175) );
  XOR2X1 U731 ( .A(n17), .B(n995), .Y(n1177) );
  XOR2X1 U732 ( .A(n936), .B(n937), .Y(n935) );
  XOR2X1 U733 ( .A(n938), .B(n806), .Y(n937) );
  XOR2X1 U734 ( .A(n55), .B(n939), .Y(n936) );
  XOR2X1 U735 ( .A(n134), .B(n756), .Y(n938) );
  XOR2X1 U736 ( .A(n408), .B(n409), .Y(n407) );
  XOR2X1 U737 ( .A(n299), .B(n410), .Y(n409) );
  XOR2X1 U738 ( .A(n282), .B(n411), .Y(n408) );
  XOR2X1 U739 ( .A(round_key[108]), .B(new_block[4]), .Y(n411) );
  XOR2X1 U740 ( .A(n1198), .B(n1199), .Y(n1197) );
  XOR2X1 U741 ( .A(n1200), .B(n1045), .Y(n1199) );
  XOR2X1 U742 ( .A(n82), .B(n1201), .Y(n1198) );
  XOR2X1 U743 ( .A(n20), .B(n1022), .Y(n1200) );
  XOR2X1 U744 ( .A(n718), .B(n719), .Y(n717) );
  XOR2X1 U745 ( .A(n720), .B(n565), .Y(n719) );
  XOR2X1 U746 ( .A(n146), .B(n721), .Y(n718) );
  XOR2X1 U747 ( .A(n90), .B(n542), .Y(n720) );
  XOR2X1 U748 ( .A(n849), .B(n850), .Y(n848) );
  XOR2X1 U749 ( .A(n851), .B(n790), .Y(n850) );
  XOR2X1 U750 ( .A(n28), .B(n852), .Y(n849) );
  XOR2X1 U751 ( .A(n138), .B(n740), .Y(n851) );
  XOR2X1 U752 ( .A(n571), .B(n572), .Y(n570) );
  XOR2X1 U753 ( .A(new_block[13]), .B(n506), .Y(n572) );
  XOR2X1 U754 ( .A(new_block[53]), .B(n573), .Y(n571) );
  XOR2X1 U755 ( .A(round_key[86]), .B(new_block[94]), .Y(n573) );
  XOR2X1 U756 ( .A(n471), .B(n472), .Y(n470) );
  XOR2X1 U757 ( .A(n473), .B(n333), .Y(n472) );
  XOR2X1 U758 ( .A(n42), .B(n474), .Y(n471) );
  XOR2X1 U759 ( .A(n120), .B(n289), .Y(n473) );
  XOR2X1 U760 ( .A(n479), .B(n480), .Y(n478) );
  XOR2X1 U761 ( .A(new_block[121]), .B(n300), .Y(n480) );
  XOR2X1 U762 ( .A(new_block[1]), .B(n481), .Y(n479) );
  XOR2X1 U763 ( .A(round_key[98]), .B(new_block[42]), .Y(n481) );
  XOR2X1 U764 ( .A(round_key[126]), .B(new_block[86]), .Y(n271) );
  XOR2X1 U765 ( .A(round_key[125]), .B(new_block[85]), .Y(n279) );
  XOR2X1 U766 ( .A(round_key[122]), .B(new_block[82]), .Y(n306) );
  XOR2X1 U767 ( .A(round_key[120]), .B(new_block[80]), .Y(n323) );
  XOR2X1 U768 ( .A(round_key[127]), .B(new_block[7]), .Y(n263) );
  XOR2X1 U769 ( .A(round_key[63]), .B(new_block[71]), .Y(n737) );
  XOR2X1 U770 ( .A(n875), .B(n876), .Y(n874) );
  XOR2X1 U771 ( .A(n748), .B(n765), .Y(n876) );
  XOR2X1 U772 ( .A(round_key[45]), .B(new_block[69]), .Y(n875) );
  XOR2X1 U773 ( .A(n402), .B(n403), .Y(n401) );
  XOR2X1 U774 ( .A(n274), .B(n291), .Y(n403) );
  XOR2X1 U775 ( .A(round_key[109]), .B(new_block[5]), .Y(n402) );
  XOR2X1 U776 ( .A(n396), .B(n397), .Y(n395) );
  XOR2X1 U777 ( .A(n265), .B(n281), .Y(n397) );
  XOR2X1 U778 ( .A(round_key[110]), .B(new_block[6]), .Y(n396) );
  XOR2X1 U779 ( .A(n869), .B(n870), .Y(n868) );
  XOR2X1 U780 ( .A(n739), .B(n755), .Y(n870) );
  XOR2X1 U781 ( .A(round_key[46]), .B(new_block[70]), .Y(n869) );
  XOR2X1 U782 ( .A(n655), .B(n656), .Y(n654) );
  XOR2X1 U783 ( .A(n533), .B(n549), .Y(n656) );
  XOR2X1 U784 ( .A(round_key[74]), .B(new_block[98]), .Y(n655) );
  XOR2X1 U785 ( .A(n390), .B(n391), .Y(n389) );
  XOR2X1 U786 ( .A(n273), .B(n333), .Y(n391) );
  XOR2X1 U787 ( .A(round_key[111]), .B(new_block[87]), .Y(n390) );
  XOR2X1 U788 ( .A(n896), .B(n897), .Y(n895) );
  XOR2X1 U789 ( .A(n774), .B(n790), .Y(n897) );
  XOR2X1 U790 ( .A(round_key[42]), .B(new_block[66]), .Y(n896) );
  XOR2X1 U791 ( .A(n1206), .B(n1207), .Y(n1205) );
  XOR2X1 U792 ( .A(n1030), .B(n1045), .Y(n1207) );
  XOR2X1 U793 ( .A(round_key[0]), .B(new_block[72]), .Y(n1206) );
  XOR2X1 U794 ( .A(round_key[62]), .B(new_block[22]), .Y(n745) );
  XOR2X1 U795 ( .A(round_key[31]), .B(new_block[39]), .Y(n976) );
  XOR2X1 U796 ( .A(round_key[94]), .B(new_block[54]), .Y(n504) );
  XOR2X1 U797 ( .A(n1108), .B(n1109), .Y(n1107) );
  XOR2X1 U798 ( .A(n978), .B(n994), .Y(n1109) );
  XOR2X1 U799 ( .A(round_key[14]), .B(new_block[38]), .Y(n1108) );
  XOR2X1 U800 ( .A(n863), .B(n864), .Y(n862) );
  XOR2X1 U801 ( .A(n747), .B(n806), .Y(n864) );
  XOR2X1 U802 ( .A(round_key[47]), .B(new_block[23]), .Y(n863) );
  XOR2X1 U803 ( .A(n622), .B(n623), .Y(n621) );
  XOR2X1 U804 ( .A(n506), .B(n565), .Y(n623) );
  XOR2X1 U805 ( .A(round_key[79]), .B(new_block[55]), .Y(n622) );
  XOR2X1 U806 ( .A(n726), .B(n727), .Y(n725) );
  XOR2X1 U807 ( .A(n550), .B(n565), .Y(n727) );
  XOR2X1 U808 ( .A(round_key[64]), .B(new_block[8]), .Y(n726) );
  XOR2X1 U809 ( .A(round_key[29]), .B(new_block[117]), .Y(n992) );
  XOR2X1 U810 ( .A(round_key[61]), .B(new_block[21]), .Y(n753) );
  XOR2X1 U811 ( .A(round_key[30]), .B(new_block[118]), .Y(n984) );
  XOR2X1 U812 ( .A(round_key[93]), .B(new_block[53]), .Y(n512) );
  XOR2X1 U813 ( .A(round_key[95]), .B(new_block[103]), .Y(n496) );
  XOR2X1 U814 ( .A(n628), .B(n629), .Y(n627) );
  XOR2X1 U815 ( .A(n498), .B(n514), .Y(n629) );
  XOR2X1 U816 ( .A(round_key[78]), .B(new_block[102]), .Y(n628) );
  XOR2X1 U817 ( .A(n634), .B(n635), .Y(n633) );
  XOR2X1 U818 ( .A(n507), .B(n524), .Y(n635) );
  XOR2X1 U819 ( .A(round_key[77]), .B(new_block[101]), .Y(n634) );
  XOR2X1 U820 ( .A(n1114), .B(n1115), .Y(n1113) );
  XOR2X1 U821 ( .A(n987), .B(n1004), .Y(n1115) );
  XOR2X1 U822 ( .A(round_key[13]), .B(new_block[37]), .Y(n1114) );
  XOR2X1 U823 ( .A(n1102), .B(n1103), .Y(n1101) );
  XOR2X1 U824 ( .A(n986), .B(n1045), .Y(n1103) );
  XOR2X1 U825 ( .A(round_key[15]), .B(new_block[119]), .Y(n1102) );
  XOR2X1 U826 ( .A(n384), .B(n385), .Y(n383) );
  XOR2X1 U827 ( .A(n266), .B(n325), .Y(n385) );
  XOR2X1 U828 ( .A(round_key[112]), .B(new_block[120]), .Y(n384) );
  XOR2X1 U829 ( .A(round_key[26]), .B(new_block[114]), .Y(n1019) );
  XOR2X1 U830 ( .A(round_key[56]), .B(new_block[16]), .Y(n797) );
  XOR2X1 U831 ( .A(round_key[58]), .B(new_block[18]), .Y(n780) );
  XOR2X1 U832 ( .A(round_key[24]), .B(new_block[112]), .Y(n1036) );
  XOR2X1 U833 ( .A(round_key[90]), .B(new_block[50]), .Y(n539) );
  XOR2X1 U834 ( .A(round_key[88]), .B(new_block[48]), .Y(n556) );
  XOR2X1 U835 ( .A(n967), .B(n968), .Y(n966) );
  XOR2X1 U836 ( .A(n791), .B(n806), .Y(n968) );
  XOR2X1 U837 ( .A(round_key[32]), .B(new_block[104]), .Y(n967) );
  XOR2X1 U838 ( .A(n331), .B(n332), .Y(n330) );
  XOR2X1 U839 ( .A(new_block[46]), .B(n333), .Y(n332) );
  XOR2X1 U840 ( .A(new_block[47]), .B(n334), .Y(n331) );
  XOR2X1 U841 ( .A(round_key[119]), .B(new_block[86]), .Y(n334) );
  XOR2X1 U842 ( .A(n563), .B(n564), .Y(n562) );
  XOR2X1 U843 ( .A(new_block[14]), .B(n565), .Y(n564) );
  XOR2X1 U844 ( .A(new_block[15]), .B(n566), .Y(n563) );
  XOR2X1 U845 ( .A(round_key[87]), .B(new_block[54]), .Y(n566) );
  XOR2X1 U846 ( .A(n804), .B(n805), .Y(n803) );
  XOR2X1 U847 ( .A(new_block[110]), .B(n806), .Y(n805) );
  XOR2X1 U848 ( .A(new_block[111]), .B(n807), .Y(n804) );
  XOR2X1 U849 ( .A(round_key[55]), .B(new_block[22]), .Y(n807) );
  XOR2X1 U850 ( .A(n1043), .B(n1044), .Y(n1042) );
  XOR2X1 U851 ( .A(new_block[118]), .B(n1045), .Y(n1044) );
  XOR2X1 U852 ( .A(new_block[78]), .B(n1046), .Y(n1043) );
  XOR2X1 U853 ( .A(round_key[23]), .B(new_block[79]), .Y(n1046) );
  XOR2X1 U854 ( .A(n1183), .B(n1184), .Y(n1182) );
  XOR2X1 U855 ( .A(n1185), .B(n1045), .Y(n1184) );
  XOR2X1 U856 ( .A(n80), .B(n1186), .Y(n1183) );
  XOR2X1 U857 ( .A(n18), .B(n1002), .Y(n1185) );
  XOR2X1 U858 ( .A(n944), .B(n945), .Y(n943) );
  XOR2X1 U859 ( .A(n946), .B(n806), .Y(n945) );
  XOR2X1 U860 ( .A(n56), .B(n947), .Y(n944) );
  XOR2X1 U861 ( .A(n135), .B(n763), .Y(n946) );
  XOR2X1 U862 ( .A(n703), .B(n704), .Y(n702) );
  XOR2X1 U863 ( .A(n705), .B(n565), .Y(n704) );
  XOR2X1 U864 ( .A(n88), .B(n706), .Y(n703) );
  XOR2X1 U865 ( .A(n33), .B(n522), .Y(n705) );
  XOR2X1 U866 ( .A(n1213), .B(n1214), .Y(n1212) );
  XOR2X1 U867 ( .A(n317), .B(n333), .Y(n1214) );
  XOR2X1 U868 ( .A(round_key[96]), .B(new_block[40]), .Y(n1213) );
  XOR2X1 U869 ( .A(n695), .B(n696), .Y(n694) );
  XOR2X1 U870 ( .A(n697), .B(n565), .Y(n696) );
  XOR2X1 U871 ( .A(n87), .B(n698), .Y(n695) );
  XOR2X1 U872 ( .A(n32), .B(n515), .Y(n697) );
  XOR2X1 U873 ( .A(n463), .B(n464), .Y(n462) );
  XOR2X1 U874 ( .A(n465), .B(n333), .Y(n464) );
  XOR2X1 U875 ( .A(n41), .B(n466), .Y(n463) );
  XOR2X1 U876 ( .A(n119), .B(n282), .Y(n465) );
  XOR2X1 U877 ( .A(n959), .B(n960), .Y(n958) );
  XOR2X1 U878 ( .A(n961), .B(n806), .Y(n960) );
  XOR2X1 U879 ( .A(n58), .B(n962), .Y(n959) );
  XOR2X1 U880 ( .A(n137), .B(n783), .Y(n961) );
  XOR2X1 U881 ( .A(n486), .B(n487), .Y(n485) );
  XOR2X1 U882 ( .A(n488), .B(n333), .Y(n487) );
  XOR2X1 U883 ( .A(n122), .B(n489), .Y(n486) );
  XOR2X1 U884 ( .A(n44), .B(n309), .Y(n488) );
  XOR2X1 U885 ( .A(n674), .B(n675), .Y(n673) );
  XOR2X1 U886 ( .A(new_block[102]), .B(n499), .Y(n675) );
  XOR2X1 U887 ( .A(new_block[94]), .B(n676), .Y(n674) );
  XOR2X1 U888 ( .A(round_key[71]), .B(new_block[95]), .Y(n676) );
  XOR2X1 U889 ( .A(n915), .B(n916), .Y(n914) );
  XOR2X1 U890 ( .A(new_block[62]), .B(n740), .Y(n916) );
  XOR2X1 U891 ( .A(new_block[63]), .B(n917), .Y(n915) );
  XOR2X1 U892 ( .A(round_key[39]), .B(new_block[70]), .Y(n917) );
  XOR2X1 U893 ( .A(n1154), .B(n1155), .Y(n1153) );
  XOR2X1 U894 ( .A(new_block[30]), .B(n979), .Y(n1155) );
  XOR2X1 U895 ( .A(new_block[31]), .B(n1156), .Y(n1154) );
  XOR2X1 U896 ( .A(round_key[7]), .B(new_block[38]), .Y(n1156) );
  XOR2X1 U897 ( .A(n442), .B(n443), .Y(n441) );
  XOR2X1 U898 ( .A(new_block[126]), .B(n266), .Y(n443) );
  XOR2X1 U899 ( .A(new_block[127]), .B(n444), .Y(n442) );
  XOR2X1 U900 ( .A(round_key[103]), .B(new_block[6]), .Y(n444) );
  XOR2X1 U901 ( .A(n1128), .B(n1129), .Y(n1127) );
  XOR2X1 U902 ( .A(n1021), .B(n1122), .Y(n1129) );
  XOR2X1 U903 ( .A(n1002), .B(n1130), .Y(n1128) );
  XOR2X1 U904 ( .A(round_key[11]), .B(new_block[35]), .Y(n1130) );
  XOR2X1 U905 ( .A(n889), .B(n890), .Y(n888) );
  XOR2X1 U906 ( .A(n782), .B(n883), .Y(n890) );
  XOR2X1 U907 ( .A(n763), .B(n891), .Y(n889) );
  XOR2X1 U908 ( .A(round_key[43]), .B(new_block[67]), .Y(n891) );
  XOR2X1 U909 ( .A(n416), .B(n417), .Y(n415) );
  XOR2X1 U910 ( .A(n308), .B(n410), .Y(n417) );
  XOR2X1 U911 ( .A(n289), .B(n418), .Y(n416) );
  XOR2X1 U912 ( .A(round_key[107]), .B(new_block[3]), .Y(n418) );
  XOR2X1 U913 ( .A(n648), .B(n649), .Y(n647) );
  XOR2X1 U914 ( .A(n541), .B(n642), .Y(n649) );
  XOR2X1 U915 ( .A(n522), .B(n650), .Y(n648) );
  XOR2X1 U916 ( .A(round_key[75]), .B(new_block[99]), .Y(n650) );
  XOR2X1 U917 ( .A(n1120), .B(n1121), .Y(n1119) );
  XOR2X1 U918 ( .A(n1012), .B(n1122), .Y(n1121) );
  XOR2X1 U919 ( .A(n995), .B(n1123), .Y(n1120) );
  XOR2X1 U920 ( .A(round_key[12]), .B(new_block[36]), .Y(n1123) );
  XOR2X1 U921 ( .A(n1141), .B(n1142), .Y(n1140) );
  XOR2X1 U922 ( .A(n1038), .B(n1122), .Y(n1142) );
  XOR2X1 U923 ( .A(n1022), .B(n1143), .Y(n1141) );
  XOR2X1 U924 ( .A(round_key[9]), .B(new_block[33]), .Y(n1143) );
  XOR2X1 U925 ( .A(n429), .B(n430), .Y(n428) );
  XOR2X1 U926 ( .A(n325), .B(n410), .Y(n430) );
  XOR2X1 U927 ( .A(n309), .B(n431), .Y(n429) );
  XOR2X1 U928 ( .A(round_key[105]), .B(new_block[1]), .Y(n431) );
  XOR2X1 U929 ( .A(n640), .B(n641), .Y(n639) );
  XOR2X1 U930 ( .A(n532), .B(n642), .Y(n641) );
  XOR2X1 U931 ( .A(n515), .B(n643), .Y(n640) );
  XOR2X1 U932 ( .A(round_key[76]), .B(new_block[100]), .Y(n643) );
  XOR2X1 U933 ( .A(n661), .B(n662), .Y(n660) );
  XOR2X1 U934 ( .A(n558), .B(n642), .Y(n662) );
  XOR2X1 U935 ( .A(n542), .B(n663), .Y(n661) );
  XOR2X1 U936 ( .A(round_key[73]), .B(new_block[97]), .Y(n663) );
  XOR2X1 U937 ( .A(n520), .B(n521), .Y(n517) );
  XOR2X1 U938 ( .A(n522), .B(n523), .Y(n521) );
  XOR2X1 U939 ( .A(n524), .B(n525), .Y(n520) );
  XOR2X1 U940 ( .A(round_key[92]), .B(new_block[52]), .Y(n525) );
  XOR2X1 U941 ( .A(n1000), .B(n1001), .Y(n997) );
  XOR2X1 U942 ( .A(n1002), .B(n1003), .Y(n1001) );
  XOR2X1 U943 ( .A(n1004), .B(n1005), .Y(n1000) );
  XOR2X1 U944 ( .A(round_key[28]), .B(new_block[116]), .Y(n1005) );
  XOR2X1 U945 ( .A(n761), .B(n762), .Y(n758) );
  XOR2X1 U946 ( .A(n763), .B(n764), .Y(n762) );
  XOR2X1 U947 ( .A(n765), .B(n766), .Y(n761) );
  XOR2X1 U948 ( .A(round_key[60]), .B(new_block[20]), .Y(n766) );
  XOR2X1 U949 ( .A(n771), .B(n772), .Y(n768) );
  XOR2X1 U950 ( .A(n773), .B(n774), .Y(n772) );
  XOR2X1 U951 ( .A(n764), .B(n775), .Y(n771) );
  XOR2X1 U952 ( .A(round_key[59]), .B(new_block[19]), .Y(n775) );
  XOR2X1 U953 ( .A(n1010), .B(n1011), .Y(n1007) );
  XOR2X1 U954 ( .A(n1012), .B(n1013), .Y(n1011) );
  XOR2X1 U955 ( .A(n1003), .B(n1014), .Y(n1010) );
  XOR2X1 U956 ( .A(round_key[27]), .B(new_block[115]), .Y(n1014) );
  XOR2X1 U957 ( .A(n530), .B(n531), .Y(n527) );
  XOR2X1 U958 ( .A(n532), .B(n533), .Y(n531) );
  XOR2X1 U959 ( .A(n523), .B(n534), .Y(n530) );
  XOR2X1 U960 ( .A(round_key[91]), .B(new_block[51]), .Y(n534) );
  XOR2X1 U961 ( .A(n1027), .B(n1028), .Y(n1024) );
  XOR2X1 U962 ( .A(n1029), .B(n1030), .Y(n1028) );
  XOR2X1 U963 ( .A(n1003), .B(n1031), .Y(n1027) );
  XOR2X1 U964 ( .A(round_key[25]), .B(new_block[113]), .Y(n1031) );
  XOR2X1 U965 ( .A(n788), .B(n789), .Y(n785) );
  XOR2X1 U966 ( .A(n790), .B(n791), .Y(n789) );
  XOR2X1 U967 ( .A(n764), .B(n792), .Y(n788) );
  XOR2X1 U968 ( .A(round_key[57]), .B(new_block[17]), .Y(n792) );
  XOR2X1 U969 ( .A(n547), .B(n548), .Y(n544) );
  XOR2X1 U970 ( .A(n549), .B(n550), .Y(n548) );
  XOR2X1 U971 ( .A(n523), .B(n551), .Y(n547) );
  XOR2X1 U972 ( .A(round_key[89]), .B(new_block[49]), .Y(n551) );
  XOR2X1 U973 ( .A(n353), .B(n354), .Y(n352) );
  XOR2X1 U974 ( .A(n355), .B(n291), .Y(n354) );
  XOR2X1 U975 ( .A(n71), .B(n356), .Y(n353) );
  XOR2X1 U976 ( .A(n118), .B(n266), .Y(n355) );
  XOR2X1 U977 ( .A(n826), .B(n827), .Y(n825) );
  XOR2X1 U978 ( .A(n828), .B(n765), .Y(n827) );
  XOR2X1 U979 ( .A(n25), .B(n829), .Y(n826) );
  XOR2X1 U980 ( .A(n135), .B(n740), .Y(n828) );
  XOR2X1 U981 ( .A(n1065), .B(n1066), .Y(n1064) );
  XOR2X1 U982 ( .A(n1067), .B(n1004), .Y(n1066) );
  XOR2X1 U983 ( .A(n16), .B(n1068), .Y(n1065) );
  XOR2X1 U984 ( .A(n127), .B(n979), .Y(n1067) );
  XOR2X1 U985 ( .A(n608), .B(n609), .Y(n607) );
  XOR2X1 U986 ( .A(n610), .B(n549), .Y(n609) );
  XOR2X1 U987 ( .A(n89), .B(n611), .Y(n608) );
  XOR2X1 U988 ( .A(n66), .B(n499), .Y(n610) );
  XOR2X1 U989 ( .A(n1088), .B(n1089), .Y(n1087) );
  XOR2X1 U990 ( .A(n1090), .B(n1029), .Y(n1089) );
  XOR2X1 U991 ( .A(n19), .B(n1091), .Y(n1088) );
  XOR2X1 U992 ( .A(n130), .B(n979), .Y(n1090) );
  XOR2X1 U993 ( .A(n857), .B(n858), .Y(n856) );
  XOR2X1 U994 ( .A(n740), .B(n799), .Y(n858) );
  XOR2X1 U995 ( .A(round_key[48]), .B(new_block[56]), .Y(n857) );
  XOR2X1 U996 ( .A(n819), .B(n820), .Y(n818) );
  XOR2X1 U997 ( .A(new_block[108]), .B(n755), .Y(n820) );
  XOR2X1 U998 ( .A(new_block[20]), .B(n821), .Y(n819) );
  XOR2X1 U999 ( .A(round_key[53]), .B(new_block[61]), .Y(n821) );
  XOR2X1 U1000 ( .A(n1096), .B(n1097), .Y(n1095) );
  XOR2X1 U1001 ( .A(n979), .B(n1038), .Y(n1097) );
  XOR2X1 U1002 ( .A(round_key[16]), .B(new_block[24]), .Y(n1096) );
  XOR2X1 U1003 ( .A(n346), .B(n347), .Y(n345) );
  XOR2X1 U1004 ( .A(new_block[125]), .B(n281), .Y(n347) );
  XOR2X1 U1005 ( .A(new_block[44]), .B(n348), .Y(n346) );
  XOR2X1 U1006 ( .A(round_key[117]), .B(new_block[84]), .Y(n348) );
  XOR2X1 U1007 ( .A(n1135), .B(n1136), .Y(n1134) );
  XOR2X1 U1008 ( .A(n1013), .B(n1029), .Y(n1136) );
  XOR2X1 U1009 ( .A(round_key[10]), .B(new_block[34]), .Y(n1135) );
  XOR2X1 U1010 ( .A(n688), .B(n689), .Y(n687) );
  XOR2X1 U1011 ( .A(new_block[100]), .B(n507), .Y(n689) );
  XOR2X1 U1012 ( .A(new_block[13]), .B(n690), .Y(n688) );
  XOR2X1 U1013 ( .A(round_key[69]), .B(new_block[92]), .Y(n690) );
  XOR2X1 U1014 ( .A(n456), .B(n457), .Y(n455) );
  XOR2X1 U1015 ( .A(new_block[124]), .B(n274), .Y(n457) );
  XOR2X1 U1016 ( .A(new_block[45]), .B(n458), .Y(n456) );
  XOR2X1 U1017 ( .A(round_key[101]), .B(new_block[4]), .Y(n458) );
  XOR2X1 U1018 ( .A(n376), .B(n377), .Y(n375) );
  XOR2X1 U1019 ( .A(n378), .B(n316), .Y(n377) );
  XOR2X1 U1020 ( .A(n74), .B(n379), .Y(n376) );
  XOR2X1 U1021 ( .A(n121), .B(n266), .Y(n378) );
  XOR2X1 U1022 ( .A(n929), .B(n930), .Y(n928) );
  XOR2X1 U1023 ( .A(new_block[109]), .B(n748), .Y(n930) );
  XOR2X1 U1024 ( .A(new_block[60]), .B(n931), .Y(n929) );
  XOR2X1 U1025 ( .A(round_key[37]), .B(new_block[68]), .Y(n931) );
  XOR2X1 U1026 ( .A(n423), .B(n424), .Y(n422) );
  XOR2X1 U1027 ( .A(n300), .B(n316), .Y(n424) );
  XOR2X1 U1028 ( .A(round_key[106]), .B(new_block[2]), .Y(n423) );
  XOR2X1 U1029 ( .A(n578), .B(n579), .Y(n577) );
  XOR2X1 U1030 ( .A(new_block[12]), .B(n514), .Y(n579) );
  XOR2X1 U1031 ( .A(new_block[52]), .B(n580), .Y(n578) );
  XOR2X1 U1032 ( .A(round_key[85]), .B(new_block[93]), .Y(n580) );
  XOR2X1 U1033 ( .A(n1168), .B(n1169), .Y(n1167) );
  XOR2X1 U1034 ( .A(new_block[28]), .B(n987), .Y(n1169) );
  XOR2X1 U1035 ( .A(new_block[36]), .B(n1170), .Y(n1168) );
  XOR2X1 U1036 ( .A(round_key[5]), .B(new_block[77]), .Y(n1170) );
  XOR2X1 U1037 ( .A(n616), .B(n617), .Y(n615) );
  XOR2X1 U1038 ( .A(n499), .B(n558), .Y(n617) );
  XOR2X1 U1039 ( .A(round_key[80]), .B(new_block[88]), .Y(n616) );
  XOR2X1 U1040 ( .A(n952), .B(n953), .Y(n951) );
  XOR2X1 U1041 ( .A(new_block[106]), .B(n774), .Y(n953) );
  XOR2X1 U1042 ( .A(new_block[57]), .B(n954), .Y(n952) );
  XOR2X1 U1043 ( .A(round_key[34]), .B(new_block[65]), .Y(n954) );
  XOR2X1 U1044 ( .A(n585), .B(n586), .Y(n584) );
  XOR2X1 U1045 ( .A(n587), .B(n524), .Y(n586) );
  XOR2X1 U1046 ( .A(n63), .B(n588), .Y(n585) );
  XOR2X1 U1047 ( .A(n33), .B(n499), .Y(n587) );
  XOR2X1 U1048 ( .A(n1191), .B(n1192), .Y(n1190) );
  XOR2X1 U1049 ( .A(new_block[25]), .B(n1013), .Y(n1192) );
  XOR2X1 U1050 ( .A(new_block[33]), .B(n1193), .Y(n1191) );
  XOR2X1 U1051 ( .A(round_key[2]), .B(new_block[74]), .Y(n1193) );
  XOR2X1 U1052 ( .A(n711), .B(n712), .Y(n710) );
  XOR2X1 U1053 ( .A(new_block[10]), .B(n533), .Y(n712) );
  XOR2X1 U1054 ( .A(new_block[89]), .B(n713), .Y(n711) );
  XOR2X1 U1055 ( .A(round_key[66]), .B(new_block[97]), .Y(n713) );
  XOR2X1 U1056 ( .A(n593), .B(n594), .Y(n592) );
  XOR2X1 U1057 ( .A(n595), .B(n532), .Y(n594) );
  XOR2X1 U1058 ( .A(n64), .B(n596), .Y(n593) );
  XOR2X1 U1059 ( .A(n34), .B(n499), .Y(n595) );
  XOR2X1 U1060 ( .A(n834), .B(n835), .Y(n833) );
  XOR2X1 U1061 ( .A(n836), .B(n773), .Y(n835) );
  XOR2X1 U1062 ( .A(n26), .B(n837), .Y(n834) );
  XOR2X1 U1063 ( .A(n136), .B(n740), .Y(n836) );
  XOR2X1 U1064 ( .A(n1073), .B(n1074), .Y(n1072) );
  XOR2X1 U1065 ( .A(n1075), .B(n1012), .Y(n1074) );
  XOR2X1 U1066 ( .A(n17), .B(n1076), .Y(n1073) );
  XOR2X1 U1067 ( .A(n128), .B(n979), .Y(n1075) );
  XOR2X1 U1068 ( .A(n601), .B(n602), .Y(n600) );
  XOR2X1 U1069 ( .A(new_block[49]), .B(n541), .Y(n602) );
  XOR2X1 U1070 ( .A(new_block[90]), .B(n603), .Y(n601) );
  XOR2X1 U1071 ( .A(round_key[82]), .B(new_block[9]), .Y(n603) );
  XOR2X1 U1072 ( .A(n842), .B(n843), .Y(n841) );
  XOR2X1 U1073 ( .A(new_block[105]), .B(n782), .Y(n843) );
  XOR2X1 U1074 ( .A(new_block[17]), .B(n844), .Y(n842) );
  XOR2X1 U1075 ( .A(round_key[50]), .B(new_block[58]), .Y(n844) );
  XOR2X1 U1076 ( .A(n1081), .B(n1082), .Y(n1080) );
  XOR2X1 U1077 ( .A(new_block[113]), .B(n1021), .Y(n1082) );
  XOR2X1 U1078 ( .A(new_block[26]), .B(n1083), .Y(n1081) );
  XOR2X1 U1079 ( .A(round_key[18]), .B(new_block[73]), .Y(n1083) );
  XOR2X1 U1080 ( .A(n339), .B(n340), .Y(n338) );
  XOR2X1 U1081 ( .A(new_block[126]), .B(n273), .Y(n340) );
  XOR2X1 U1082 ( .A(new_block[45]), .B(n341), .Y(n339) );
  XOR2X1 U1083 ( .A(round_key[118]), .B(new_block[85]), .Y(n341) );
  XOR2X1 U1084 ( .A(n812), .B(n813), .Y(n811) );
  XOR2X1 U1085 ( .A(new_block[109]), .B(n747), .Y(n813) );
  XOR2X1 U1086 ( .A(new_block[21]), .B(n814), .Y(n812) );
  XOR2X1 U1087 ( .A(round_key[54]), .B(new_block[62]), .Y(n814) );
  XOR2X1 U1088 ( .A(n1051), .B(n1052), .Y(n1050) );
  XOR2X1 U1089 ( .A(new_block[117]), .B(n986), .Y(n1052) );
  XOR2X1 U1090 ( .A(new_block[30]), .B(n1053), .Y(n1051) );
  XOR2X1 U1091 ( .A(round_key[22]), .B(new_block[77]), .Y(n1053) );
  XOR2X1 U1092 ( .A(n361), .B(n362), .Y(n360) );
  XOR2X1 U1093 ( .A(n363), .B(n299), .Y(n362) );
  XOR2X1 U1094 ( .A(n72), .B(n364), .Y(n361) );
  XOR2X1 U1095 ( .A(n119), .B(n266), .Y(n363) );
  XOR2X1 U1096 ( .A(n369), .B(n370), .Y(n368) );
  XOR2X1 U1097 ( .A(new_block[122]), .B(n308), .Y(n370) );
  XOR2X1 U1098 ( .A(new_block[41]), .B(n371), .Y(n369) );
  XOR2X1 U1099 ( .A(round_key[114]), .B(new_block[81]), .Y(n371) );
  XOR2X1 U1100 ( .A(n449), .B(n450), .Y(n448) );
  XOR2X1 U1101 ( .A(new_block[125]), .B(n265), .Y(n450) );
  XOR2X1 U1102 ( .A(new_block[46]), .B(n451), .Y(n449) );
  XOR2X1 U1103 ( .A(round_key[102]), .B(new_block[5]), .Y(n451) );
  XOR2X1 U1104 ( .A(n681), .B(n682), .Y(n680) );
  XOR2X1 U1105 ( .A(new_block[101]), .B(n498), .Y(n682) );
  XOR2X1 U1106 ( .A(new_block[14]), .B(n683), .Y(n681) );
  XOR2X1 U1107 ( .A(round_key[70]), .B(new_block[93]), .Y(n683) );
  XOR2X1 U1108 ( .A(n1161), .B(n1162), .Y(n1160) );
  XOR2X1 U1109 ( .A(new_block[29]), .B(n978), .Y(n1162) );
  XOR2X1 U1110 ( .A(new_block[37]), .B(n1163), .Y(n1161) );
  XOR2X1 U1111 ( .A(round_key[6]), .B(new_block[78]), .Y(n1163) );
  OAI22XL U1112 ( .A0(block[93]), .A1(n177), .B0(new_block[93]), .B1(n162), 
        .Y(n511) );
  OAI22XL U1113 ( .A0(block[92]), .A1(n177), .B0(new_block[92]), .B1(n162), 
        .Y(n519) );
  OAI22XL U1114 ( .A0(block[95]), .A1(n187), .B0(new_block[95]), .B1(n161), 
        .Y(n495) );
  OAI22XL U1115 ( .A0(block[62]), .A1(n190), .B0(new_block[62]), .B1(n162), 
        .Y(n744) );
  OAI22XL U1116 ( .A0(block[61]), .A1(n189), .B0(new_block[61]), .B1(n163), 
        .Y(n752) );
  OAI22XL U1117 ( .A0(block[60]), .A1(n191), .B0(new_block[60]), .B1(n163), 
        .Y(n760) );
  OAI22XL U1118 ( .A0(block[57]), .A1(n189), .B0(new_block[57]), .B1(n163), 
        .Y(n787) );
  OAI22XL U1119 ( .A0(block[94]), .A1(n187), .B0(new_block[94]), .B1(n161), 
        .Y(n503) );
  OAI22XL U1120 ( .A0(block[29]), .A1(n188), .B0(new_block[29]), .B1(n163), 
        .Y(n991) );
  OAI22XL U1121 ( .A0(block[31]), .A1(n190), .B0(new_block[31]), .B1(n163), 
        .Y(n975) );
  OAI22XL U1122 ( .A0(block[30]), .A1(n189), .B0(new_block[30]), .B1(n163), 
        .Y(n983) );
  OAI22XL U1123 ( .A0(block[63]), .A1(n191), .B0(new_block[63]), .B1(n162), 
        .Y(n736) );
  OAI22XL U1124 ( .A0(block[126]), .A1(n190), .B0(new_block[126]), .B1(n161), 
        .Y(n270) );
  OAI22XL U1125 ( .A0(block[125]), .A1(n189), .B0(new_block[125]), .B1(n161), 
        .Y(n278) );
  OAI22XL U1126 ( .A0(block[127]), .A1(n189), .B0(new_block[127]), .B1(n162), 
        .Y(n261) );
  OAI22XL U1127 ( .A0(n52), .A1(n159), .B0(n176), .B1(n1458), .Y(n743) );
  INVX1 U1128 ( .A(block[62]), .Y(n1458) );
  OAI22XL U1129 ( .A0(n15), .A1(n158), .B0(n192), .B1(n1455), .Y(n990) );
  INVX1 U1130 ( .A(block[29]), .Y(n1455) );
  OAI22XL U1131 ( .A0(n18), .A1(n158), .B0(n176), .B1(n1443), .Y(n1017) );
  INVX1 U1132 ( .A(block[26]), .Y(n1443) );
  OAI22XL U1133 ( .A0(n58), .A1(n158), .B0(n192), .B1(n1438), .Y(n795) );
  INVX1 U1134 ( .A(block[56]), .Y(n1438) );
  OAI22XL U1135 ( .A0(n53), .A1(n160), .B0(n176), .B1(n1454), .Y(n751) );
  INVX1 U1136 ( .A(block[61]), .Y(n1454) );
  OAI22XL U1137 ( .A0(n56), .A1(n159), .B0(n187), .B1(n1442), .Y(n778) );
  INVX1 U1138 ( .A(block[58]), .Y(n1442) );
  OAI22XL U1139 ( .A0(n20), .A1(n158), .B0(n176), .B1(n1439), .Y(n1034) );
  INVX1 U1140 ( .A(block[24]), .Y(n1439) );
  OAI22XL U1141 ( .A0(n13), .A1(n159), .B0(n192), .B1(n1463), .Y(n974) );
  INVX1 U1142 ( .A(block[31]), .Y(n1463) );
  OAI22XL U1143 ( .A0(n14), .A1(n159), .B0(n176), .B1(n1459), .Y(n982) );
  INVX1 U1144 ( .A(block[30]), .Y(n1459) );
  OAI22XL U1145 ( .A0(n116), .A1(n158), .B0(n187), .B1(n1456), .Y(n269) );
  INVX1 U1146 ( .A(block[126]), .Y(n1456) );
  OAI22XL U1147 ( .A0(n117), .A1(n158), .B0(n190), .B1(n1452), .Y(n277) );
  INVX1 U1148 ( .A(block[125]), .Y(n1452) );
  OAI22XL U1149 ( .A0(n120), .A1(n159), .B0(n189), .B1(n1440), .Y(n304) );
  INVX1 U1150 ( .A(block[122]), .Y(n1440) );
  OAI22XL U1151 ( .A0(n122), .A1(n160), .B0(n191), .B1(n1436), .Y(n321) );
  INVX1 U1152 ( .A(block[120]), .Y(n1436) );
  OAI22XL U1153 ( .A0(n115), .A1(n158), .B0(n188), .B1(n1460), .Y(n260) );
  INVX1 U1154 ( .A(block[127]), .Y(n1460) );
  OAI22XL U1155 ( .A0(n84), .A1(n160), .B0(n176), .B1(n1457), .Y(n502) );
  INVX1 U1156 ( .A(block[94]), .Y(n1457) );
  OAI22XL U1157 ( .A0(n85), .A1(n161), .B0(n176), .B1(n1453), .Y(n510) );
  INVX1 U1158 ( .A(block[93]), .Y(n1453) );
  OAI22XL U1159 ( .A0(n88), .A1(n160), .B0(n176), .B1(n1441), .Y(n537) );
  INVX1 U1160 ( .A(block[90]), .Y(n1441) );
  OAI22XL U1161 ( .A0(n90), .A1(n160), .B0(n192), .B1(n1437), .Y(n554) );
  INVX1 U1162 ( .A(block[88]), .Y(n1437) );
  OAI22XL U1163 ( .A0(n83), .A1(n159), .B0(n190), .B1(n1461), .Y(n494) );
  INVX1 U1164 ( .A(block[95]), .Y(n1461) );
  OAI22XL U1165 ( .A0(n51), .A1(n160), .B0(n262), .B1(n1462), .Y(n735) );
  INVX1 U1166 ( .A(block[63]), .Y(n1462) );
  OAI22XL U1167 ( .A0(block[56]), .A1(n190), .B0(new_block[56]), .B1(n163), 
        .Y(n796) );
  OAI22XL U1168 ( .A0(block[59]), .A1(n191), .B0(new_block[59]), .B1(n163), 
        .Y(n770) );
  OAI22XL U1169 ( .A0(block[58]), .A1(n188), .B0(new_block[58]), .B1(n163), 
        .Y(n779) );
  OAI22XL U1170 ( .A0(block[24]), .A1(n187), .B0(new_block[24]), .B1(n164), 
        .Y(n1035) );
  OAI22XL U1171 ( .A0(block[91]), .A1(n177), .B0(new_block[91]), .B1(n162), 
        .Y(n529) );
  OAI22XL U1172 ( .A0(block[88]), .A1(n177), .B0(new_block[88]), .B1(n162), 
        .Y(n555) );
  OAI22XL U1173 ( .A0(block[28]), .A1(n188), .B0(new_block[28]), .B1(n163), 
        .Y(n999) );
  OAI22XL U1174 ( .A0(block[26]), .A1(n177), .B0(new_block[26]), .B1(n164), 
        .Y(n1018) );
  OAI22XL U1175 ( .A0(block[25]), .A1(n177), .B0(new_block[25]), .B1(n164), 
        .Y(n1026) );
  OAI22XL U1176 ( .A0(block[120]), .A1(n191), .B0(new_block[120]), .B1(n162), 
        .Y(n322) );
  OAI22XL U1177 ( .A0(block[90]), .A1(n177), .B0(new_block[90]), .B1(n162), 
        .Y(n538) );
  OAI22XL U1178 ( .A0(block[89]), .A1(n177), .B0(new_block[89]), .B1(n162), 
        .Y(n546) );
  OAI22XL U1179 ( .A0(block[27]), .A1(n177), .B0(new_block[27]), .B1(n164), 
        .Y(n1009) );
  OAI22XL U1180 ( .A0(block[124]), .A1(n191), .B0(new_block[124]), .B1(n161), 
        .Y(n286) );
  OAI22XL U1181 ( .A0(block[123]), .A1(n177), .B0(new_block[123]), .B1(n161), 
        .Y(n296) );
  OAI22XL U1182 ( .A0(block[122]), .A1(n188), .B0(new_block[122]), .B1(n161), 
        .Y(n305) );
  OAI22XL U1183 ( .A0(block[121]), .A1(n190), .B0(new_block[121]), .B1(n161), 
        .Y(n313) );
  XOR2X1 U1184 ( .A(new_block[103]), .B(new_block[95]), .Y(n565) );
  XOR2X1 U1185 ( .A(new_block[63]), .B(new_block[71]), .Y(n806) );
  XOR2X1 U1186 ( .A(new_block[127]), .B(new_block[7]), .Y(n333) );
  XOR2X1 U1187 ( .A(new_block[31]), .B(new_block[39]), .Y(n1045) );
  XOR2X1 U1188 ( .A(new_block[119]), .B(new_block[79]), .Y(n979) );
  XOR2X1 U1189 ( .A(new_block[47]), .B(new_block[87]), .Y(n266) );
  XOR2X1 U1190 ( .A(new_block[15]), .B(new_block[55]), .Y(n499) );
  XOR2X1 U1191 ( .A(new_block[111]), .B(new_block[23]), .Y(n740) );
  XOR2X1 U1192 ( .A(new_block[123]), .B(new_block[83]), .Y(n289) );
  XOR2X1 U1193 ( .A(n909), .B(n910), .Y(n908) );
  XOR2X1 U1194 ( .A(n791), .B(n883), .Y(n910) );
  XOR2X1 U1195 ( .A(round_key[40]), .B(new_block[64]), .Y(n909) );
  XOR2X1 U1196 ( .A(n668), .B(n669), .Y(n667) );
  XOR2X1 U1197 ( .A(n550), .B(n642), .Y(n669) );
  XOR2X1 U1198 ( .A(round_key[72]), .B(new_block[96]), .Y(n668) );
  XOR2X1 U1199 ( .A(n1148), .B(n1149), .Y(n1147) );
  XOR2X1 U1200 ( .A(n1030), .B(n1122), .Y(n1149) );
  XOR2X1 U1201 ( .A(round_key[8]), .B(new_block[32]), .Y(n1148) );
  XOR2X1 U1202 ( .A(n436), .B(n437), .Y(n435) );
  XOR2X1 U1203 ( .A(n317), .B(n410), .Y(n437) );
  XOR2X1 U1204 ( .A(round_key[104]), .B(new_block[0]), .Y(n436) );
  XOR2X1 U1205 ( .A(round_key[96]), .B(new_block[0]), .Y(n1211) );
  OAI2BB1X1 U1206 ( .A0N(ready), .A1N(n1220), .B0(n164), .Y(n1361) );
  XOR2X1 U1207 ( .A(new_block[39]), .B(new_block[79]), .Y(n1122) );
  XOR2X1 U1208 ( .A(new_block[111]), .B(new_block[71]), .Y(n883) );
  XOR2X1 U1209 ( .A(new_block[47]), .B(new_block[7]), .Y(n410) );
  XOR2X1 U1210 ( .A(new_block[103]), .B(new_block[15]), .Y(n642) );
  XOR2X1 U1211 ( .A(new_block[55]), .B(new_block[95]), .Y(n523) );
  XOR2X1 U1212 ( .A(new_block[127]), .B(new_block[87]), .Y(n290) );
  XOR2X1 U1213 ( .A(new_block[23]), .B(new_block[63]), .Y(n764) );
  XOR2X1 U1214 ( .A(new_block[119]), .B(new_block[31]), .Y(n1003) );
  XOR2X1 U1215 ( .A(new_block[52]), .B(new_block[92]), .Y(n515) );
  XOR2X1 U1216 ( .A(new_block[53]), .B(new_block[93]), .Y(n507) );
  XOR2X1 U1217 ( .A(new_block[97]), .B(new_block[9]), .Y(n549) );
  XOR2X1 U1218 ( .A(new_block[108]), .B(new_block[68]), .Y(n765) );
  XOR2X1 U1219 ( .A(new_block[124]), .B(new_block[84]), .Y(n282) );
  XOR2X1 U1220 ( .A(new_block[44]), .B(new_block[4]), .Y(n291) );
  XOR2X1 U1221 ( .A(new_block[121]), .B(new_block[81]), .Y(n309) );
  XOR2X1 U1222 ( .A(new_block[45]), .B(new_block[5]), .Y(n281) );
  XOR2X1 U1223 ( .A(new_block[109]), .B(new_block[69]), .Y(n755) );
  XOR2X1 U1224 ( .A(new_block[37]), .B(new_block[77]), .Y(n994) );
  XOR2X1 U1225 ( .A(new_block[36]), .B(new_block[76]), .Y(n1004) );
  XOR2X1 U1226 ( .A(new_block[33]), .B(new_block[73]), .Y(n1029) );
  XOR2X1 U1227 ( .A(new_block[32]), .B(new_block[72]), .Y(n1038) );
  XOR2X1 U1228 ( .A(new_block[125]), .B(new_block[85]), .Y(n274) );
  XOR2X1 U1229 ( .A(new_block[105]), .B(new_block[65]), .Y(n790) );
  XOR2X1 U1230 ( .A(new_block[122]), .B(new_block[82]), .Y(n300) );
  XOR2X1 U1231 ( .A(new_block[104]), .B(new_block[64]), .Y(n799) );
  XOR2X1 U1232 ( .A(new_block[20]), .B(new_block[60]), .Y(n756) );
  XOR2X1 U1233 ( .A(new_block[17]), .B(new_block[57]), .Y(n783) );
  XOR2X1 U1234 ( .A(new_block[21]), .B(new_block[61]), .Y(n748) );
  XOR2X1 U1235 ( .A(new_block[1]), .B(new_block[41]), .Y(n316) );
  XOR2X1 U1236 ( .A(new_block[117]), .B(new_block[29]), .Y(n987) );
  XOR2X1 U1237 ( .A(new_block[101]), .B(new_block[13]), .Y(n514) );
  XOR2X1 U1238 ( .A(new_block[18]), .B(new_block[58]), .Y(n774) );
  XOR2X1 U1239 ( .A(new_block[8]), .B(new_block[96]), .Y(n558) );
  XOR2X1 U1240 ( .A(new_block[0]), .B(new_block[40]), .Y(n325) );
  XOR2X1 U1241 ( .A(new_block[116]), .B(new_block[28]), .Y(n995) );
  XOR2X1 U1242 ( .A(new_block[49]), .B(new_block[89]), .Y(n542) );
  XOR2X1 U1243 ( .A(new_block[113]), .B(new_block[25]), .Y(n1022) );
  XOR2X1 U1244 ( .A(new_block[114]), .B(new_block[26]), .Y(n1013) );
  XOR2X1 U1245 ( .A(new_block[50]), .B(new_block[90]), .Y(n533) );
  XOR2X1 U1246 ( .A(new_block[100]), .B(new_block[12]), .Y(n524) );
  XOR2X1 U1247 ( .A(new_block[11]), .B(new_block[99]), .Y(n532) );
  XOR2X1 U1248 ( .A(new_block[35]), .B(new_block[75]), .Y(n1012) );
  XOR2X1 U1249 ( .A(new_block[10]), .B(new_block[98]), .Y(n541) );
  XOR2X1 U1250 ( .A(new_block[34]), .B(new_block[74]), .Y(n1021) );
  XOR2X1 U1251 ( .A(new_block[110]), .B(new_block[70]), .Y(n747) );
  XOR2X1 U1252 ( .A(new_block[46]), .B(new_block[6]), .Y(n273) );
  XOR2X1 U1253 ( .A(new_block[126]), .B(new_block[86]), .Y(n265) );
  XOR2X1 U1254 ( .A(new_block[107]), .B(new_block[67]), .Y(n773) );
  XOR2X1 U1255 ( .A(new_block[106]), .B(new_block[66]), .Y(n782) );
  XOR2X1 U1256 ( .A(new_block[120]), .B(new_block[80]), .Y(n317) );
  XOR2X1 U1257 ( .A(new_block[22]), .B(new_block[62]), .Y(n739) );
  XOR2X1 U1258 ( .A(new_block[54]), .B(new_block[94]), .Y(n498) );
  XOR2X1 U1259 ( .A(new_block[38]), .B(new_block[78]), .Y(n986) );
  XOR2X1 U1260 ( .A(new_block[118]), .B(new_block[30]), .Y(n978) );
  XOR2X1 U1261 ( .A(new_block[102]), .B(new_block[14]), .Y(n506) );
  XOR2X1 U1262 ( .A(new_block[19]), .B(new_block[59]), .Y(n763) );
  XOR2X1 U1263 ( .A(new_block[51]), .B(new_block[91]), .Y(n522) );
  XOR2X1 U1264 ( .A(new_block[112]), .B(new_block[24]), .Y(n1030) );
  XOR2X1 U1265 ( .A(new_block[16]), .B(new_block[56]), .Y(n791) );
  XOR2X1 U1266 ( .A(new_block[48]), .B(new_block[88]), .Y(n550) );
  XOR2X1 U1267 ( .A(new_block[3]), .B(new_block[43]), .Y(n299) );
  XOR2X1 U1268 ( .A(new_block[2]), .B(new_block[42]), .Y(n308) );
  XOR2X1 U1269 ( .A(new_block[115]), .B(new_block[27]), .Y(n1002) );
  OAI22XL U1270 ( .A0(n48), .A1(n1227), .B0(round[0]), .B1(n1431), .Y(n1365)
         );
  NAND3X1 U1271 ( .A(n12), .B(n11), .C(next), .Y(n1220) );
  NAND4X1 U1272 ( .A(round[2]), .B(n1223), .C(round[1]), .D(n45), .Y(n1222) );
  NAND2X1 U1273 ( .A(n11), .B(next), .Y(n1232) );
  OA21XL U1274 ( .A0(round[1]), .A1(n1431), .B0(n1226), .Y(n1225) );
  OA21XL U1275 ( .A0(round[0]), .A1(n1431), .B0(n1227), .Y(n1226) );
  OAI211X1 U1276 ( .A0(enc_ctrl_we), .A1(n12), .B0(n1220), .C0(n1228), .Y(
        n1366) );
  OAI211X1 U1277 ( .A0(enc_ctrl_we), .A1(n11), .B0(n1429), .C0(n1228), .Y(
        n1367) );
  OAI22XL U1278 ( .A0(n50), .A1(n1230), .B0(sword_ctr_reg[0]), .B1(n1219), .Y(
        n1369) );
  OAI22XL U1279 ( .A0(n49), .A1(n1230), .B0(n1231), .B1(n1219), .Y(n1368) );
  NOR2X1 U1280 ( .A(n730), .B(n969), .Y(n1231) );
  INVX1 U1281 ( .A(block[28]), .Y(n1451) );
  INVX1 U1282 ( .A(block[27]), .Y(n1447) );
  INVX1 U1283 ( .A(block[25]), .Y(n1434) );
  INVX1 U1284 ( .A(block[60]), .Y(n1450) );
  INVX1 U1285 ( .A(block[59]), .Y(n1446) );
  INVX1 U1286 ( .A(block[57]), .Y(n1432) );
  INVX1 U1287 ( .A(block[124]), .Y(n1448) );
  INVX1 U1288 ( .A(block[123]), .Y(n1444) );
  INVX1 U1289 ( .A(block[121]), .Y(n1433) );
  INVX1 U1290 ( .A(block[92]), .Y(n1449) );
  INVX1 U1291 ( .A(block[91]), .Y(n1445) );
  INVX1 U1292 ( .A(block[89]), .Y(n1435) );
  OAI221XL U1293 ( .A0(n482), .A1(n183), .B0(n145), .B1(n207), .C0(n483), .Y(
        n1263) );
  OAI221XL U1294 ( .A0(n714), .A1(n179), .B0(n113), .B1(n155), .C0(n715), .Y(
        n1294) );
  OAI221XL U1295 ( .A0(n955), .A1(n182), .B0(n81), .B1(n152), .C0(n956), .Y(
        n1326) );
  OAI221XL U1296 ( .A0(n1194), .A1(n186), .B0(n43), .B1(n149), .C0(n1195), .Y(
        n1358) );
  OAI221XL U1297 ( .A0(n404), .A1(n184), .B0(n134), .B1(n1), .C0(n405), .Y(
        n1252) );
  OAI221XL U1298 ( .A0(n636), .A1(n180), .B0(n102), .B1(n156), .C0(n637), .Y(
        n1283) );
  OAI221XL U1299 ( .A0(n877), .A1(n178), .B0(n70), .B1(n153), .C0(n878), .Y(
        n1315) );
  OAI221XL U1300 ( .A0(n1116), .A1(n185), .B0(n32), .B1(n150), .C0(n1117), .Y(
        n1347) );
  OAI221XL U1301 ( .A0(n432), .A1(n183), .B0(n138), .B1(n207), .C0(n433), .Y(
        n1256) );
  OAI221XL U1302 ( .A0(n664), .A1(n180), .B0(n106), .B1(n155), .C0(n665), .Y(
        n1287) );
  OAI221XL U1303 ( .A0(n905), .A1(n179), .B0(n74), .B1(n152), .C0(n906), .Y(
        n1319) );
  OAI221XL U1304 ( .A0(n1144), .A1(n186), .B0(n36), .B1(n149), .C0(n1145), .Y(
        n1351) );
  OAI221XL U1305 ( .A0(n459), .A1(n183), .B0(n142), .B1(n207), .C0(n460), .Y(
        n1260) );
  OAI221XL U1306 ( .A0(n691), .A1(n179), .B0(n110), .B1(n155), .C0(n692), .Y(
        n1291) );
  OAI221XL U1307 ( .A0(n932), .A1(n181), .B0(n78), .B1(n152), .C0(n933), .Y(
        n1323) );
  OAI221XL U1308 ( .A0(n1171), .A1(n186), .B0(n40), .B1(n149), .C0(n1172), .Y(
        n1355) );
  OR2X1 U1309 ( .A(n1221), .B(n40), .Y(n3) );
  NAND2X1 U1310 ( .A(n729), .B(n210), .Y(n732) );
  OA22XL U1311 ( .A0(n222), .A1(n83), .B0(n211), .B1(n51), .Y(n230) );
  OA22XL U1312 ( .A0(n222), .A1(n84), .B0(n211), .B1(n52), .Y(n231) );
  OA22XL U1313 ( .A0(n215), .A1(n85), .B0(n211), .B1(n53), .Y(n233) );
  OA22XL U1314 ( .A0(n215), .A1(n87), .B0(n211), .B1(n55), .Y(n235) );
  OA22XL U1315 ( .A0(n215), .A1(n86), .B0(n211), .B1(n54), .Y(n234) );
  OAI221XL U1316 ( .A0(n219), .A1(n21), .B0(n216), .B1(n123), .C0(n239), .Y(
        sboxw[23]) );
  OAI221XL U1317 ( .A0(n219), .A1(n22), .B0(n216), .B1(n124), .C0(n240), .Y(
        sboxw[22]) );
  OAI221XL U1318 ( .A0(n1224), .A1(n23), .B0(n216), .B1(n125), .C0(n241), .Y(
        sboxw[21]) );
  OAI221XL U1319 ( .A0(n1224), .A1(n26), .B0(n216), .B1(n128), .C0(n245), .Y(
        sboxw[18]) );
  OAI221XL U1320 ( .A0(n219), .A1(n18), .B0(n216), .B1(n120), .C0(n236), .Y(
        sboxw[26]) );
  OAI221XL U1321 ( .A0(n1224), .A1(n24), .B0(n216), .B1(n126), .C0(n242), .Y(
        sboxw[20]) );
  OAI221XL U1322 ( .A0(n1224), .A1(n25), .B0(n216), .B1(n127), .C0(n244), .Y(
        sboxw[19]) );
  OA22XL U1323 ( .A0(n215), .A1(n107), .B0(n212), .B1(n75), .Y(n225) );
  OA22XL U1324 ( .A0(n214), .A1(n91), .B0(n223), .B1(n59), .Y(n239) );
  OA22XL U1325 ( .A0(n214), .A1(n92), .B0(n223), .B1(n60), .Y(n240) );
  OA22XL U1326 ( .A0(n214), .A1(n93), .B0(n212), .B1(n61), .Y(n241) );
  OA22XL U1327 ( .A0(n214), .A1(n96), .B0(n212), .B1(n64), .Y(n245) );
  OA22XL U1328 ( .A0(n214), .A1(n88), .B0(n223), .B1(n56), .Y(n236) );
  OA22XL U1329 ( .A0(n214), .A1(n94), .B0(n212), .B1(n62), .Y(n242) );
  OA22XL U1330 ( .A0(n214), .A1(n95), .B0(n212), .B1(n63), .Y(n244) );
  OA22XL U1331 ( .A0(n214), .A1(n90), .B0(n212), .B1(n58), .Y(n238) );
  OA22XL U1332 ( .A0(n214), .A1(n89), .B0(n212), .B1(n57), .Y(n237) );
  AOI222XL U1333 ( .A0(new_sboxw[6]), .A1(n1426), .B0(n171), .B1(n447), .C0(
        n201), .C1(n448), .Y(n446) );
  AOI222XL U1334 ( .A0(n5), .A1(new_sboxw[6]), .B0(n168), .B1(n679), .C0(n198), 
        .C1(n680), .Y(n678) );
  AOI222XL U1335 ( .A0(n147), .A1(new_sboxw[6]), .B0(n174), .B1(n920), .C0(
        n201), .C1(n921), .Y(n919) );
  AOI222XL U1336 ( .A0(n9), .A1(new_sboxw[6]), .B0(n173), .B1(n1159), .C0(n194), .C1(n1160), .Y(n1158) );
  OA22XL U1337 ( .A0(n213), .A1(n98), .B0(n210), .B1(n66), .Y(n247) );
  OA22XL U1338 ( .A0(n213), .A1(n97), .B0(n210), .B1(n65), .Y(n246) );
  AOI222XL U1339 ( .A0(new_sboxw[1]), .A1(n8), .B0(n170), .B1(n484), .C0(n195), 
        .C1(n485), .Y(n483) );
  AOI222XL U1340 ( .A0(n5), .A1(new_sboxw[1]), .B0(n168), .B1(n716), .C0(n198), 
        .C1(n717), .Y(n715) );
  AOI222XL U1341 ( .A0(n147), .A1(new_sboxw[1]), .B0(n175), .B1(n957), .C0(
        n201), .C1(n958), .Y(n956) );
  AOI222XL U1342 ( .A0(n9), .A1(new_sboxw[1]), .B0(n328), .B1(n1196), .C0(n193), .C1(n1197), .Y(n1195) );
  AOI222XL U1343 ( .A0(new_sboxw[8]), .A1(n8), .B0(n171), .B1(n434), .C0(n205), 
        .C1(n435), .Y(n433) );
  AOI222XL U1344 ( .A0(n5), .A1(new_sboxw[8]), .B0(n169), .B1(n666), .C0(n197), 
        .C1(n667), .Y(n665) );
  AOI222XL U1345 ( .A0(n147), .A1(new_sboxw[8]), .B0(n175), .B1(n907), .C0(
        n201), .C1(n908), .Y(n906) );
  AOI222XL U1346 ( .A0(n9), .A1(new_sboxw[8]), .B0(n174), .B1(n1146), .C0(n195), .C1(n1147), .Y(n1145) );
  OAI22XL U1347 ( .A0(n1226), .A1(n47), .B0(round[1]), .B1(n1430), .Y(n1364)
         );
  OAI32XL U1348 ( .A0(n1430), .A1(round[2]), .A2(n47), .B0(n1225), .B1(n46), 
        .Y(n1363) );
  AOI222XL U1349 ( .A0(new_sboxw[9]), .A1(n8), .B0(n171), .B1(n427), .C0(n204), 
        .C1(n428), .Y(n426) );
  AOI222XL U1350 ( .A0(n5), .A1(new_sboxw[9]), .B0(n169), .B1(n659), .C0(n197), 
        .C1(n660), .Y(n658) );
  AOI222XL U1351 ( .A0(n147), .A1(new_sboxw[9]), .B0(n165), .B1(n900), .C0(
        n200), .C1(n901), .Y(n899) );
  AOI222XL U1352 ( .A0(n9), .A1(new_sboxw[9]), .B0(n174), .B1(n1139), .C0(n195), .C1(n1140), .Y(n1138) );
  NOR2BXL U1353 ( .AN(n1217), .B(n1218), .Y(n328) );
  AOI222XL U1354 ( .A0(new_sboxw[4]), .A1(n8), .B0(n171), .B1(n461), .C0(n195), 
        .C1(n462), .Y(n460) );
  AOI222XL U1355 ( .A0(n5), .A1(new_sboxw[4]), .B0(n168), .B1(n693), .C0(n198), 
        .C1(n694), .Y(n692) );
  AOI222XL U1356 ( .A0(n147), .A1(new_sboxw[4]), .B0(n175), .B1(n934), .C0(
        n201), .C1(n935), .Y(n933) );
  AOI222XL U1357 ( .A0(n9), .A1(new_sboxw[4]), .B0(n166), .B1(n1173), .C0(n193), .C1(n1174), .Y(n1172) );
  NAND2X1 U1358 ( .A(n1216), .B(n1215), .Y(n262) );
  AOI222XL U1359 ( .A0(new_sboxw[12]), .A1(n7), .B0(n171), .B1(n406), .C0(n203), .C1(n407), .Y(n405) );
  AOI222XL U1360 ( .A0(n6), .A1(new_sboxw[12]), .B0(n169), .B1(n638), .C0(n197), .C1(n639), .Y(n637) );
  AOI222XL U1361 ( .A0(n148), .A1(new_sboxw[12]), .B0(n167), .B1(n879), .C0(
        n200), .C1(n880), .Y(n878) );
  AOI222XL U1362 ( .A0(n10), .A1(new_sboxw[12]), .B0(n173), .B1(n1118), .C0(
        n195), .C1(n1119), .Y(n1117) );
endmodule


module aes_inv_sbox ( sword, new_sword );
  input [31:0] sword;
  output [31:0] new_sword;
  wire   n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n363, n579, n906, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548;

  INVX1 U1 ( .A(n903), .Y(n1446) );
  INVX1 U2 ( .A(n142), .Y(n1497) );
  INVX1 U3 ( .A(n360), .Y(n1521) );
  INVX1 U4 ( .A(n1443), .Y(n36) );
  INVX1 U5 ( .A(n1494), .Y(n62) );
  INVX1 U6 ( .A(n1518), .Y(n73) );
  NOR2X1 U7 ( .A(n1506), .B(n64), .Y(n720) );
  NOR2X1 U8 ( .A(n1455), .B(n38), .Y(n1016) );
  NOR2X1 U9 ( .A(n1534), .B(n75), .Y(n473) );
  INVX1 U10 ( .A(n1220), .Y(n201) );
  INVX1 U11 ( .A(n3), .Y(n123) );
  INVX1 U12 ( .A(n1), .Y(n133) );
  INVX1 U13 ( .A(n2), .Y(n106) );
  OAI222XL U14 ( .A0(n130), .A1(n1439), .B0(n125), .B1(n35), .C0(n101), .C1(
        n42), .Y(n1059) );
  OAI222XL U15 ( .A0(n407), .A1(n1514), .B0(n108), .B1(n72), .C0(n93), .C1(n79), .Y(n516) );
  OAI222XL U16 ( .A0(n623), .A1(n1490), .B0(n135), .B1(n61), .C0(n105), .C1(
        n68), .Y(n763) );
  NOR2X1 U17 ( .A(n203), .B(n227), .Y(n1220) );
  NOR2X1 U18 ( .A(n226), .B(n205), .Y(n269) );
  NOR2X1 U19 ( .A(n224), .B(n205), .Y(n294) );
  NOR2X1 U20 ( .A(n64), .B(n1504), .Y(n649) );
  NOR2X1 U21 ( .A(n38), .B(n1453), .Y(n976) );
  NOR2X1 U22 ( .A(n75), .B(n1532), .Y(n433) );
  OR2X1 U23 ( .A(n58), .B(n103), .Y(n1) );
  OR2X1 U24 ( .A(n45), .B(n91), .Y(n2) );
  NOR2X1 U25 ( .A(n38), .B(n1457), .Y(n918) );
  NOR2X1 U26 ( .A(n64), .B(n1507), .Y(n591) );
  NOR2X1 U27 ( .A(n75), .B(n1535), .Y(n375) );
  INVX1 U28 ( .A(n284), .Y(n212) );
  INVX1 U29 ( .A(n424), .Y(n1520) );
  INVX1 U30 ( .A(n967), .Y(n1445) );
  INVX1 U31 ( .A(n640), .Y(n1496) );
  OR2X1 U32 ( .A(n32), .B(n99), .Y(n3) );
  OAI22XL U33 ( .A0(sword[18]), .A1(n28), .B0(n38), .B1(n1425), .Y(n1020) );
  OAI22XL U34 ( .A0(sword[2]), .A1(n11), .B0(n75), .B1(n179), .Y(n477) );
  OAI22XL U35 ( .A0(sword[26]), .A1(n54), .B0(n64), .B1(n1476), .Y(n724) );
  NOR2X1 U36 ( .A(n227), .B(sword[11]), .Y(n289) );
  OAI22XL U37 ( .A0(n205), .A1(n147), .B0(sword[10]), .B1(n143), .Y(n1322) );
  NOR2X1 U38 ( .A(n225), .B(sword[10]), .Y(n284) );
  NOR2X1 U39 ( .A(n70), .B(sword[26]), .Y(n640) );
  NOR2X1 U40 ( .A(n44), .B(sword[18]), .Y(n967) );
  NOR2X1 U41 ( .A(n81), .B(sword[2]), .Y(n424) );
  NOR2X1 U42 ( .A(n220), .B(sword[12]), .Y(n1248) );
  NOR2X1 U43 ( .A(n203), .B(sword[12]), .Y(n1210) );
  INVX1 U44 ( .A(sword[10]), .Y(n205) );
  NOR2X1 U45 ( .A(n1492), .B(sword[28]), .Y(n574) );
  NOR2X1 U46 ( .A(n1441), .B(sword[20]), .Y(n901) );
  NOR2X1 U47 ( .A(n1516), .B(sword[4]), .Y(n358) );
  NOR2X1 U48 ( .A(n1535), .B(sword[3]), .Y(n400) );
  NOR2X1 U49 ( .A(n1457), .B(sword[19]), .Y(n943) );
  NOR2X1 U50 ( .A(n1507), .B(sword[27]), .Y(n616) );
  INVX1 U51 ( .A(sword[20]), .Y(n1457) );
  INVX1 U52 ( .A(sword[4]), .Y(n1535) );
  INVX1 U53 ( .A(sword[28]), .Y(n1507) );
  INVX1 U54 ( .A(sword[12]), .Y(n227) );
  NOR2X1 U55 ( .A(n1453), .B(sword[20]), .Y(n908) );
  NOR2X1 U56 ( .A(n1504), .B(sword[28]), .Y(n581) );
  NOR2X1 U57 ( .A(n1532), .B(sword[4]), .Y(n365) );
  NOR2X1 U58 ( .A(n224), .B(sword[12]), .Y(n307) );
  NOR2X1 U59 ( .A(n205), .B(sword[11]), .Y(n1227) );
  NOR2X1 U60 ( .A(n39), .B(sword[19]), .Y(n978) );
  NOR2X1 U61 ( .A(n76), .B(sword[3]), .Y(n435) );
  NOR2X1 U62 ( .A(n65), .B(sword[27]), .Y(n651) );
  INVX1 U63 ( .A(sword[14]), .Y(n233) );
  INVX1 U64 ( .A(sword[22]), .Y(n1463) );
  INVX1 U65 ( .A(sword[6]), .Y(n1541) );
  INVX1 U66 ( .A(sword[30]), .Y(n1527) );
  BUFX2 U67 ( .A(n1421), .Y(n22) );
  BUFX2 U68 ( .A(n1472), .Y(n47) );
  BUFX2 U69 ( .A(n175), .Y(n4) );
  INVX1 U70 ( .A(n268), .Y(n82) );
  INVX1 U71 ( .A(n129), .Y(n25) );
  INVX1 U72 ( .A(n112), .Y(n8) );
  INVX1 U73 ( .A(n139), .Y(n51) );
  INVX1 U74 ( .A(n122), .Y(n83) );
  INVX1 U75 ( .A(n399), .Y(n183) );
  INVX1 U76 ( .A(n942), .Y(n1429) );
  INVX1 U77 ( .A(n615), .Y(n1480) );
  INVX1 U78 ( .A(n890), .Y(n26) );
  INVX1 U79 ( .A(n139), .Y(n52) );
  INVX1 U80 ( .A(n112), .Y(n9) );
  INVX1 U81 ( .A(n506), .Y(n180) );
  INVX1 U82 ( .A(n1049), .Y(n1426) );
  INVX1 U83 ( .A(n753), .Y(n1477) );
  BUFX2 U84 ( .A(n1544), .Y(n84) );
  BUFX2 U85 ( .A(n1472), .Y(n48) );
  BUFX2 U86 ( .A(n175), .Y(n5) );
  BUFX2 U87 ( .A(n1421), .Y(n21) );
  BUFX2 U88 ( .A(n1544), .Y(n85) );
  NOR2X1 U89 ( .A(n11), .B(n74), .Y(n399) );
  NOR2X1 U90 ( .A(n29), .B(n37), .Y(n942) );
  NOR2X1 U91 ( .A(n54), .B(n63), .Y(n615) );
  NAND4X1 U92 ( .A(n183), .B(n417), .C(n171), .D(n184), .Y(n412) );
  NAND4X1 U93 ( .A(n1429), .B(n960), .C(n1417), .D(n1430), .Y(n955) );
  NAND4X1 U94 ( .A(n1480), .B(n633), .C(n1468), .D(n1481), .Y(n628) );
  INVX1 U95 ( .A(n260), .Y(n218) );
  BUFX2 U96 ( .A(n144), .Y(n143) );
  INVX1 U97 ( .A(n1242), .Y(n196) );
  INVX1 U98 ( .A(n1318), .Y(n198) );
  INVX1 U99 ( .A(n950), .Y(n1421) );
  INVX1 U100 ( .A(n140), .Y(n1472) );
  INVX1 U101 ( .A(n113), .Y(n175) );
  NOR2X1 U102 ( .A(n74), .B(n347), .Y(n506) );
  NOR2X1 U103 ( .A(n37), .B(n129), .Y(n1049) );
  NOR2X1 U104 ( .A(n63), .B(n563), .Y(n753) );
  INVX1 U105 ( .A(n482), .Y(n181) );
  INVX1 U106 ( .A(n1025), .Y(n1427) );
  INVX1 U107 ( .A(n729), .Y(n1478) );
  INVX1 U108 ( .A(n270), .Y(n1544) );
  INVX1 U109 ( .A(n287), .Y(n217) );
  INVX1 U110 ( .A(n1019), .Y(n1432) );
  INVX1 U111 ( .A(n476), .Y(n186) );
  INVX1 U112 ( .A(n723), .Y(n1483) );
  NOR2X1 U113 ( .A(n219), .B(n122), .Y(n260) );
  NOR2X1 U114 ( .A(n16), .B(n122), .Y(n1318) );
  OAI21XL U115 ( .A0(n890), .A1(n41), .B0(n994), .Y(n1100) );
  OAI21XL U116 ( .A0(n112), .A1(n78), .B0(n451), .Y(n532) );
  OAI21XL U117 ( .A0(n139), .A1(n67), .B0(n698), .Y(n779) );
  NOR2X1 U118 ( .A(n16), .B(n1547), .Y(n1242) );
  NOR2X1 U119 ( .A(n7), .B(n77), .Y(n392) );
  NOR2X1 U120 ( .A(n24), .B(n40), .Y(n935) );
  NOR2X1 U121 ( .A(n50), .B(n66), .Y(n608) );
  BUFX2 U122 ( .A(n563), .Y(n139) );
  BUFX2 U123 ( .A(n347), .Y(n112) );
  NAND2X1 U124 ( .A(n131), .B(n25), .Y(n960) );
  NAND2X1 U125 ( .A(n114), .B(n8), .Y(n417) );
  NAND2X1 U126 ( .A(n141), .B(n51), .Y(n633) );
  NAND2X1 U127 ( .A(n131), .B(n22), .Y(n994) );
  NAND2X1 U128 ( .A(n114), .B(n4), .Y(n451) );
  NAND2X1 U129 ( .A(n141), .B(n47), .Y(n698) );
  BUFX2 U130 ( .A(n623), .Y(n140) );
  BUFX2 U131 ( .A(n407), .Y(n113) );
  BUFX2 U132 ( .A(n268), .Y(n122) );
  INVX1 U133 ( .A(n503), .Y(n184) );
  INVX1 U134 ( .A(n1046), .Y(n1430) );
  INVX1 U135 ( .A(n750), .Y(n1481) );
  INVX1 U136 ( .A(n278), .Y(n200) );
  INVX1 U137 ( .A(n454), .Y(n171) );
  INVX1 U138 ( .A(n997), .Y(n1417) );
  INVX1 U139 ( .A(n701), .Y(n1468) );
  INVX1 U140 ( .A(n116), .Y(n88) );
  INVX1 U141 ( .A(n131), .Y(n1438) );
  INVX1 U142 ( .A(n141), .Y(n1489) );
  INVX1 U143 ( .A(n114), .Y(n1513) );
  INVX1 U144 ( .A(n73), .Y(n74) );
  INVX1 U145 ( .A(n36), .Y(n37) );
  INVX1 U146 ( .A(n62), .Y(n63) );
  INVX1 U147 ( .A(n1265), .Y(n206) );
  BUFX2 U148 ( .A(n1547), .Y(n144) );
  NOR2X1 U149 ( .A(n1446), .B(n890), .Y(n1025) );
  NOR2X1 U150 ( .A(n1497), .B(n139), .Y(n729) );
  NOR2X1 U151 ( .A(n1521), .B(n112), .Y(n482) );
  NOR2X1 U152 ( .A(n1446), .B(n30), .Y(n1019) );
  NOR2X1 U153 ( .A(n1521), .B(n13), .Y(n476) );
  NOR2X1 U154 ( .A(n1497), .B(n56), .Y(n723) );
  NOR2X1 U155 ( .A(n219), .B(n84), .Y(n287) );
  NOR2X1 U156 ( .A(n40), .B(n130), .Y(n1045) );
  NOR2X1 U157 ( .A(n77), .B(n113), .Y(n502) );
  NOR2X1 U158 ( .A(n66), .B(n140), .Y(n749) );
  NOR2X1 U159 ( .A(n21), .B(n1446), .Y(n998) );
  NOR2X1 U160 ( .A(n48), .B(n1497), .Y(n702) );
  NOR2X1 U161 ( .A(n5), .B(n1521), .Y(n455) );
  BUFX2 U162 ( .A(n890), .Y(n129) );
  BUFX2 U163 ( .A(n1425), .Y(n23) );
  BUFX2 U164 ( .A(n1476), .Y(n49) );
  BUFX2 U165 ( .A(n179), .Y(n6) );
  BUFX2 U166 ( .A(n179), .Y(n7) );
  BUFX2 U167 ( .A(n1425), .Y(n24) );
  BUFX2 U168 ( .A(n1476), .Y(n50) );
  INVX1 U169 ( .A(n1368), .Y(n215) );
  INVX1 U170 ( .A(n431), .Y(n178) );
  INVX1 U171 ( .A(n974), .Y(n1424) );
  INVX1 U172 ( .A(n647), .Y(n1475) );
  BUFX2 U173 ( .A(n950), .Y(n130) );
  BUFX2 U174 ( .A(n3), .Y(n29) );
  BUFX2 U175 ( .A(n1), .Y(n55) );
  BUFX2 U176 ( .A(n2), .Y(n12) );
  INVX1 U177 ( .A(n919), .Y(n1431) );
  INVX1 U178 ( .A(n376), .Y(n185) );
  INVX1 U179 ( .A(n592), .Y(n1482) );
  BUFX2 U180 ( .A(n3), .Y(n28) );
  BUFX2 U181 ( .A(n2), .Y(n11) );
  BUFX2 U182 ( .A(n1), .Y(n54) );
  INVX1 U183 ( .A(n940), .Y(n30) );
  INVX1 U184 ( .A(n397), .Y(n13) );
  INVX1 U185 ( .A(n613), .Y(n56) );
  INVX1 U186 ( .A(n940), .Y(n31) );
  INVX1 U187 ( .A(n397), .Y(n14) );
  INVX1 U188 ( .A(n613), .Y(n57) );
  BUFX2 U189 ( .A(n270), .Y(n118) );
  INVX1 U190 ( .A(n1283), .Y(n213) );
  OAI21XL U191 ( .A0(n118), .A1(n19), .B0(n1278), .Y(n1213) );
  OAI22XL U192 ( .A0(n1547), .A1(n204), .B0(n85), .B1(n18), .Y(n321) );
  OAI22XL U193 ( .A0(n54), .A1(n1489), .B0(n48), .B1(n61), .Y(n826) );
  OAI22XL U194 ( .A0(n3), .A1(n1438), .B0(n21), .B1(n35), .Y(n1147) );
  OAI22XL U195 ( .A0(n11), .A1(n1513), .B0(n5), .B1(n72), .Y(n680) );
  NOR2X1 U196 ( .A(n201), .B(n144), .Y(n278) );
  NAND2X1 U197 ( .A(n120), .B(n144), .Y(n1253) );
  NOR2X1 U198 ( .A(n11), .B(n1514), .Y(n367) );
  NOR2X1 U199 ( .A(n28), .B(n1439), .Y(n910) );
  NOR2X1 U200 ( .A(n54), .B(n1490), .Y(n583) );
  NOR2X1 U201 ( .A(n40), .B(n27), .Y(n997) );
  NOR2X1 U202 ( .A(n77), .B(n10), .Y(n454) );
  NOR2X1 U203 ( .A(n66), .B(n53), .Y(n701) );
  NOR2X1 U204 ( .A(n1521), .B(n108), .Y(n503) );
  NOR2X1 U205 ( .A(n1446), .B(n125), .Y(n1046) );
  NOR2X1 U206 ( .A(n1497), .B(n135), .Y(n750) );
  NOR2X1 U207 ( .A(n147), .B(n207), .Y(n1265) );
  NOR2X1 U208 ( .A(n19), .B(n82), .Y(n1325) );
  NOR2X1 U209 ( .A(n33), .B(n27), .Y(n950) );
  NOR2X1 U210 ( .A(n46), .B(n10), .Y(n407) );
  NOR2X1 U211 ( .A(n145), .B(n121), .Y(n268) );
  NOR2X1 U212 ( .A(n59), .B(n53), .Y(n623) );
  NOR2X1 U213 ( .A(n123), .B(n128), .Y(n890) );
  NOR2X1 U214 ( .A(n133), .B(n138), .Y(n563) );
  NOR2X1 U215 ( .A(n106), .B(n111), .Y(n347) );
  OAI221XL U216 ( .A0(n397), .A1(n1513), .B0(n78), .B1(n4), .C0(n362), .Y(n682) );
  OAI221XL U217 ( .A0(n940), .A1(n1438), .B0(n41), .B1(n22), .C0(n905), .Y(
        n1149) );
  OAI221XL U218 ( .A0(n613), .A1(n1489), .B0(n67), .B1(n47), .C0(n578), .Y(
        n828) );
  INVX1 U219 ( .A(n148), .Y(n145) );
  NAND2X1 U220 ( .A(n117), .B(n83), .Y(n1252) );
  NAND4X1 U221 ( .A(n265), .B(n196), .C(n1252), .D(n1253), .Y(n1249) );
  OAI21XL U222 ( .A0(n129), .A1(n34), .B0(n994), .Y(n1027) );
  OAI21XL U223 ( .A0(n347), .A1(n71), .B0(n451), .Y(n484) );
  OAI21XL U224 ( .A0(n563), .A1(n60), .B0(n698), .Y(n731) );
  OAI211X1 U225 ( .A0(n1290), .A1(n83), .B0(n211), .C0(n262), .Y(n1390) );
  BUFX2 U226 ( .A(n1007), .Y(n131) );
  BUFX2 U227 ( .A(n464), .Y(n114) );
  BUFX2 U228 ( .A(n711), .Y(n141) );
  INVX1 U229 ( .A(n117), .Y(n204) );
  INVX1 U230 ( .A(n269), .Y(n15) );
  INVX1 U231 ( .A(n1016), .Y(n1443) );
  INVX1 U232 ( .A(n720), .Y(n1494) );
  INVX1 U233 ( .A(n473), .Y(n1518) );
  INVX1 U234 ( .A(n116), .Y(n1546) );
  INVX1 U235 ( .A(n885), .Y(n40) );
  INVX1 U236 ( .A(n558), .Y(n66) );
  INVX1 U237 ( .A(n342), .Y(n77) );
  INVX1 U238 ( .A(n269), .Y(n16) );
  INVX1 U239 ( .A(n558), .Y(n67) );
  INVX1 U240 ( .A(n885), .Y(n41) );
  INVX1 U241 ( .A(n342), .Y(n78) );
  INVX1 U242 ( .A(n675), .Y(n187) );
  INVX1 U243 ( .A(n1142), .Y(n1433) );
  INVX1 U244 ( .A(n821), .Y(n1484) );
  INVX1 U245 ( .A(n277), .Y(n210) );
  INVX1 U246 ( .A(n327), .Y(n208) );
  INVX1 U247 ( .A(n274), .Y(n1547) );
  INVX1 U248 ( .A(n1348), .Y(n211) );
  OAI21XL U249 ( .A0(n113), .A1(n80), .B0(n186), .Y(n346) );
  OAI21XL U250 ( .A0(n130), .A1(n43), .B0(n1432), .Y(n889) );
  OAI21XL U251 ( .A0(n140), .A1(n69), .B0(n1483), .Y(n562) );
  OAI21XL U252 ( .A0(n249), .A1(n20), .B0(n16), .Y(n1257) );
  OAI21XL U253 ( .A0(n940), .A1(n42), .B0(n37), .Y(n968) );
  OAI21XL U254 ( .A0(n397), .A1(n79), .B0(n74), .Y(n425) );
  OAI21XL U255 ( .A0(n613), .A1(n68), .B0(n63), .Y(n641) );
  NOR4X1 U256 ( .A(n1119), .B(n1024), .C(n1061), .D(n1098), .Y(n1106) );
  OAI22XL U257 ( .A0(n30), .A1(n41), .B0(n888), .B1(n1008), .Y(n1119) );
  NOR4X1 U258 ( .A(n551), .B(n481), .C(n518), .D(n530), .Y(n538) );
  OAI22XL U259 ( .A0(n13), .A1(n78), .B0(n345), .B1(n465), .Y(n551) );
  NOR2X1 U260 ( .A(n79), .B(n107), .Y(n376) );
  NOR2X1 U261 ( .A(n42), .B(n124), .Y(n919) );
  NOR2X1 U262 ( .A(n68), .B(n134), .Y(n592) );
  OAI22XL U263 ( .A0(n87), .A1(n207), .B0(n201), .B1(n83), .Y(n1281) );
  NOR2X1 U264 ( .A(n1497), .B(n53), .Y(n777) );
  NOR2X1 U265 ( .A(n1446), .B(n27), .Y(n1098) );
  NOR2X1 U266 ( .A(n1521), .B(n10), .Y(n530) );
  OAI22XL U267 ( .A0(n270), .A1(n20), .B0(n1548), .B1(n204), .Y(n1298) );
  NOR2X1 U268 ( .A(n24), .B(n43), .Y(n974) );
  NOR2X1 U269 ( .A(n7), .B(n80), .Y(n431) );
  NOR2X1 U270 ( .A(n50), .B(n69), .Y(n647) );
  NOR2X1 U271 ( .A(n20), .B(n121), .Y(n1368) );
  NOR2X1 U272 ( .A(n69), .B(n58), .Y(n765) );
  NOR2X1 U273 ( .A(n43), .B(n32), .Y(n1061) );
  NOR2X1 U274 ( .A(n80), .B(n45), .Y(n518) );
  OAI21XL U275 ( .A0(n127), .A1(n34), .B0(n1432), .Y(n1036) );
  OAI21XL U276 ( .A0(n110), .A1(n71), .B0(n186), .Y(n493) );
  OAI21XL U277 ( .A0(n137), .A1(n60), .B0(n1483), .Y(n740) );
  OAI21XL U278 ( .A0(n201), .A1(n148), .B0(n1278), .Y(n1324) );
  NOR2X1 U279 ( .A(n25), .B(n42), .Y(n1038) );
  NOR2X1 U280 ( .A(n8), .B(n79), .Y(n495) );
  NOR2X1 U281 ( .A(n51), .B(n68), .Y(n742) );
  NAND3X1 U282 ( .A(n1477), .B(n1475), .C(n854), .Y(n850) );
  AOI2BB2X1 U283 ( .B0(n135), .B1(n614), .A0N(n564), .A1N(n52), .Y(n854) );
  NAND2X1 U284 ( .A(n117), .B(n1544), .Y(n1296) );
  OA21XL U285 ( .A0(n204), .A1(n88), .B0(n19), .Y(n280) );
  OAI22XL U286 ( .A0(n84), .A1(n19), .B0(n201), .B1(n87), .Y(n1247) );
  NOR2X1 U287 ( .A(n204), .B(n86), .Y(n1232) );
  NOR2X1 U288 ( .A(n20), .B(n1546), .Y(n1283) );
  NOR4X1 U289 ( .A(n798), .B(n728), .C(n765), .D(n777), .Y(n785) );
  OAI22XL U290 ( .A0(n56), .A1(n67), .B0(n561), .B1(n712), .Y(n798) );
  NOR2X1 U291 ( .A(n23), .B(n44), .Y(n1024) );
  NOR2X1 U292 ( .A(n6), .B(n81), .Y(n481) );
  NOR2X1 U293 ( .A(n49), .B(n70), .Y(n728) );
  OAI21XL U294 ( .A0(n1007), .A1(n132), .B0(n23), .Y(n1115) );
  OAI21XL U295 ( .A0(n464), .A1(n115), .B0(n6), .Y(n547) );
  OAI21XL U296 ( .A0(n711), .A1(n576), .B0(n49), .Y(n794) );
  NOR2X1 U297 ( .A(n15), .B(n121), .Y(n282) );
  OAI21XL U298 ( .A0(n117), .A1(n120), .B0(n147), .Y(n1351) );
  NAND4BX1 U299 ( .AN(n1301), .B(n1214), .C(n1255), .D(n1296), .Y(n1365) );
  NOR2X1 U300 ( .A(n37), .B(n123), .Y(n1037) );
  NOR2X1 U301 ( .A(n63), .B(n133), .Y(n741) );
  NOR2X1 U302 ( .A(n74), .B(n106), .Y(n494) );
  NOR2X1 U303 ( .A(n1438), .B(n1428), .Y(n924) );
  NOR2X1 U304 ( .A(n1513), .B(n182), .Y(n381) );
  NOR2X1 U305 ( .A(n1489), .B(n1479), .Y(n597) );
  NOR2X1 U306 ( .A(n86), .B(n89), .Y(n270) );
  OA21XL U307 ( .A0(n14), .A1(n1513), .B0(n80), .Y(n544) );
  OA21XL U308 ( .A0(n57), .A1(n1489), .B0(n69), .Y(n791) );
  OA21XL U309 ( .A0(n31), .A1(n1438), .B0(n43), .Y(n1112) );
  OAI222XL U310 ( .A0(n32), .A1(n1438), .B0(n1443), .B1(n23), .C0(n950), .C1(
        n43), .Y(n995) );
  OAI222XL U311 ( .A0(n45), .A1(n1513), .B0(n1518), .B1(n6), .C0(n113), .C1(
        n80), .Y(n452) );
  OAI222XL U312 ( .A0(n58), .A1(n1489), .B0(n1494), .B1(n49), .C0(n140), .C1(
        n69), .Y(n699) );
  NOR2X1 U313 ( .A(n1441), .B(n33), .Y(n917) );
  NOR2X1 U314 ( .A(n1492), .B(n59), .Y(n590) );
  NOR2X1 U315 ( .A(n1516), .B(n46), .Y(n374) );
  NAND2X1 U316 ( .A(n473), .B(n182), .Y(n351) );
  NAND2X1 U317 ( .A(n1016), .B(n1428), .Y(n894) );
  NAND2X1 U318 ( .A(n720), .B(n1479), .Y(n567) );
  NAND2X1 U319 ( .A(n120), .B(n116), .Y(n1278) );
  NOR2X1 U320 ( .A(n201), .B(n1548), .Y(n1349) );
  NAND3X1 U321 ( .A(n1426), .B(n1424), .C(n1175), .Y(n1171) );
  AOI2BB2X1 U322 ( .B0(n125), .B1(n941), .A0N(n891), .A1N(n26), .Y(n1175) );
  NAND3X1 U323 ( .A(n180), .B(n178), .C(n1088), .Y(n1084) );
  AOI2BB2X1 U324 ( .B0(n108), .B1(n398), .A0N(n348), .A1N(n9), .Y(n1088) );
  INVX1 U325 ( .A(n267), .Y(n219) );
  OR4X1 U326 ( .A(n1349), .B(n282), .C(n1359), .D(n1360), .Y(n1358) );
  OAI22XL U327 ( .A0(n1547), .A1(n19), .B0(n88), .B1(n18), .Y(n1359) );
  NAND4X1 U328 ( .A(n1214), .B(n210), .C(n1296), .D(n218), .Y(n1360) );
  NOR2X1 U329 ( .A(n1548), .B(n203), .Y(n283) );
  NAND2X1 U330 ( .A(n44), .B(n1444), .Y(n1096) );
  NAND2X1 U331 ( .A(n70), .B(n1495), .Y(n775) );
  NAND2X1 U332 ( .A(n81), .B(n1519), .Y(n528) );
  INVX1 U333 ( .A(n128), .Y(n1425) );
  INVX1 U334 ( .A(n138), .Y(n1476) );
  INVX1 U335 ( .A(n111), .Y(n179) );
  NAND2X1 U336 ( .A(n66), .B(n1495), .Y(n877) );
  NAND2X1 U337 ( .A(n40), .B(n1444), .Y(n1198) );
  NAND2X1 U338 ( .A(n77), .B(n1519), .Y(n1415) );
  NAND2X1 U339 ( .A(n207), .B(n194), .Y(n332) );
  INVX1 U340 ( .A(n436), .Y(n174) );
  INVX1 U341 ( .A(n652), .Y(n1471) );
  INVX1 U342 ( .A(n979), .Y(n1420) );
  INVX1 U343 ( .A(n147), .Y(n146) );
  NAND2X1 U344 ( .A(n119), .B(n83), .Y(n1214) );
  NOR2X1 U345 ( .A(n269), .B(n1220), .Y(n1290) );
  NOR2X1 U346 ( .A(n212), .B(n116), .Y(n277) );
  NOR2X1 U347 ( .A(n1496), .B(n137), .Y(n821) );
  NOR2X1 U348 ( .A(n1445), .B(n127), .Y(n1142) );
  NOR2X1 U349 ( .A(n1520), .B(n110), .Y(n675) );
  OAI22XL U350 ( .A0(n116), .A1(n15), .B0(n222), .B1(n82), .Y(n333) );
  NOR2X1 U351 ( .A(n84), .B(n212), .Y(n327) );
  NOR2X1 U352 ( .A(n86), .B(n212), .Y(n1348) );
  NOR2X1 U353 ( .A(n1496), .B(n47), .Y(n652) );
  NOR2X1 U354 ( .A(n1445), .B(n21), .Y(n979) );
  NOR2X1 U355 ( .A(n1520), .B(n4), .Y(n436) );
  NOR2X1 U356 ( .A(n44), .B(n39), .Y(n1007) );
  NOR2X1 U357 ( .A(n81), .B(n76), .Y(n464) );
  NOR2X1 U358 ( .A(n70), .B(n65), .Y(n711) );
  OAI222XL U359 ( .A0(n127), .A1(n35), .B0(n23), .B1(n1437), .C0(n128), .C1(
        n43), .Y(n1163) );
  OAI222XL U360 ( .A0(n116), .A1(n18), .B0(n147), .B1(n192), .C0(n146), .C1(
        n19), .Y(n257) );
  OAI222XL U361 ( .A0(n137), .A1(n61), .B0(n49), .B1(n1488), .C0(n138), .C1(
        n69), .Y(n842) );
  OAI222XL U362 ( .A0(n110), .A1(n72), .B0(n6), .B1(n1512), .C0(n111), .C1(n80), .Y(n1076) );
  NOR2X1 U363 ( .A(n473), .B(n430), .Y(n465) );
  NOR2X1 U364 ( .A(n1016), .B(n973), .Y(n1008) );
  NOR2X1 U365 ( .A(n720), .B(n646), .Y(n712) );
  NAND4BX1 U366 ( .AN(n392), .B(n420), .C(n183), .D(n181), .Y(n418) );
  NAND4BX1 U367 ( .AN(n935), .B(n963), .C(n1429), .D(n1427), .Y(n961) );
  NAND4BX1 U368 ( .AN(n608), .B(n636), .C(n1480), .D(n1478), .Y(n634) );
  BUFX2 U369 ( .A(n148), .Y(n147) );
  NAND4X1 U370 ( .A(n264), .B(n262), .C(n265), .D(n266), .Y(n241) );
  AOI222XL U371 ( .A0(n267), .A1(n148), .B0(n122), .B1(n269), .C0(n118), .C1(
        n117), .Y(n266) );
  OAI21XL U372 ( .A0(n212), .A1(n88), .B0(n1253), .Y(n1205) );
  NAND4X1 U373 ( .A(n264), .B(n196), .C(n206), .D(n218), .Y(n1246) );
  OAI211X1 U374 ( .A0(n465), .A1(n9), .B0(n501), .C0(n681), .Y(n679) );
  OAI211X1 U375 ( .A0(n1008), .A1(n26), .B0(n1044), .C0(n1148), .Y(n1146) );
  OAI211X1 U376 ( .A0(n712), .A1(n52), .B0(n748), .C0(n827), .Y(n825) );
  NAND2X1 U377 ( .A(n294), .B(n82), .Y(n1217) );
  NAND2X1 U378 ( .A(n973), .B(n127), .Y(n959) );
  NAND2X1 U379 ( .A(n430), .B(n110), .Y(n416) );
  NAND2X1 U380 ( .A(n646), .B(n137), .Y(n632) );
  INVX1 U381 ( .A(n294), .Y(n203) );
  INVX1 U382 ( .A(n976), .Y(n1441) );
  INVX1 U383 ( .A(n433), .Y(n1516) );
  INVX1 U384 ( .A(n649), .Y(n1492) );
  BUFX2 U385 ( .A(n259), .Y(n117) );
  INVX1 U386 ( .A(n119), .Y(n207) );
  OAI222XL U387 ( .A0(n1506), .A1(n55), .B0(n134), .B1(n1503), .C0(n1498), 
        .C1(n52), .Y(n867) );
  OAI222XL U388 ( .A0(n1455), .A1(n29), .B0(n124), .B1(n1452), .C0(n1447), 
        .C1(n26), .Y(n1188) );
  OAI222XL U389 ( .A0(n1534), .A1(n12), .B0(n107), .B1(n1531), .C0(n1522), 
        .C1(n9), .Y(n1405) );
  BUFX2 U390 ( .A(n1545), .Y(n86) );
  AOI211X1 U391 ( .A0(n128), .A1(n132), .B0(n1100), .C0(n1048), .Y(n1099) );
  AOI211X1 U392 ( .A0(n111), .A1(n115), .B0(n532), .C0(n505), .Y(n531) );
  AOI211X1 U393 ( .A0(n138), .A1(n142), .B0(n779), .C0(n752), .Y(n778) );
  INVX1 U394 ( .A(n1248), .Y(n19) );
  INVX1 U395 ( .A(n430), .Y(n1514) );
  INVX1 U396 ( .A(n973), .Y(n1439) );
  INVX1 U397 ( .A(n646), .Y(n1490) );
  OAI211X1 U398 ( .A0(n139), .A1(n560), .B0(n568), .C0(n1497), .Y(n866) );
  OAI211X1 U399 ( .A0(n890), .A1(n887), .B0(n895), .C0(n1446), .Y(n1187) );
  OAI211X1 U400 ( .A0(n112), .A1(n344), .B0(n352), .C0(n1521), .Y(n1404) );
  BUFX2 U401 ( .A(n274), .Y(n121) );
  INVX1 U402 ( .A(n96), .Y(n89) );
  BUFX2 U403 ( .A(n888), .Y(n128) );
  BUFX2 U404 ( .A(n345), .Y(n111) );
  BUFX2 U405 ( .A(n561), .Y(n138) );
  BUFX2 U406 ( .A(n576), .Y(n142) );
  INVX1 U407 ( .A(n901), .Y(n35) );
  INVX1 U408 ( .A(n574), .Y(n61) );
  INVX1 U409 ( .A(n358), .Y(n72) );
  INVX1 U410 ( .A(n358), .Y(n71) );
  INVX1 U411 ( .A(n901), .Y(n34) );
  INVX1 U412 ( .A(n574), .Y(n60) );
  BUFX2 U413 ( .A(n1428), .Y(n27) );
  BUFX2 U414 ( .A(n182), .Y(n10) );
  BUFX2 U415 ( .A(n1479), .Y(n53) );
  INVX1 U416 ( .A(sword[25]), .Y(n58) );
  INVX1 U417 ( .A(sword[17]), .Y(n32) );
  INVX1 U418 ( .A(sword[1]), .Y(n45) );
  OAI222XL U419 ( .A0(n37), .A1(n31), .B0(n33), .B1(n999), .C0(n1451), .C1(n21), .Y(n1114) );
  OAI222XL U420 ( .A0(n74), .A1(n14), .B0(n46), .B1(n456), .C0(n1530), .C1(n5), 
        .Y(n546) );
  OAI222XL U421 ( .A0(n63), .A1(n57), .B0(n59), .B1(n703), .C0(n1502), .C1(n48), .Y(n793) );
  OAI222XL U422 ( .A0(n1546), .A1(n16), .B0(n89), .B1(n1299), .C0(n84), .C1(
        n222), .Y(n1350) );
  INVX1 U423 ( .A(n100), .Y(n33) );
  INVX1 U424 ( .A(n104), .Y(n59) );
  INVX1 U425 ( .A(n92), .Y(n46) );
  INVX1 U426 ( .A(n943), .Y(n44) );
  INVX1 U427 ( .A(n400), .Y(n81) );
  INVX1 U428 ( .A(n616), .Y(n70) );
  OA21XL U429 ( .A0(n14), .A1(n1520), .B0(n184), .Y(n362) );
  OA21XL U430 ( .A0(n31), .A1(n1445), .B0(n1430), .Y(n905) );
  OA21XL U431 ( .A0(n57), .A1(n1496), .B0(n1481), .Y(n578) );
  INVX1 U432 ( .A(n1210), .Y(n18) );
  AOI221XL U433 ( .A0(n88), .A1(n259), .B0(n118), .B1(n119), .C0(n1205), .Y(
        n1391) );
  AOI221XL U434 ( .A0(n117), .A1(n1546), .B0(n120), .B1(n121), .C0(n1375), .Y(
        n1371) );
  OAI221XL U435 ( .A0(n221), .A1(n85), .B0(n146), .B1(n1338), .C0(n1215), .Y(
        n1375) );
  INVX1 U436 ( .A(n1210), .Y(n17) );
  OAI211X1 U437 ( .A0(sword[29]), .A1(n864), .B0(n1469), .C0(n865), .Y(n858)
         );
  INVX1 U438 ( .A(n777), .Y(n1469) );
  AOI2BB2X1 U439 ( .B0(n59), .B1(n649), .A0N(n1495), .A1N(n140), .Y(n864) );
  OAI21XL U440 ( .A0(n866), .A1(n867), .B0(n164), .Y(n865) );
  OAI211X1 U441 ( .A0(sword[21]), .A1(n1185), .B0(n1418), .C0(n1186), .Y(n1179) );
  INVX1 U442 ( .A(n1098), .Y(n1418) );
  AOI2BB2X1 U443 ( .B0(n33), .B1(n976), .A0N(n1444), .A1N(n950), .Y(n1185) );
  OAI21XL U444 ( .A0(n1187), .A1(n1188), .B0(n159), .Y(n1186) );
  OAI211X1 U445 ( .A0(sword[5]), .A1(n1402), .B0(n172), .C0(n1403), .Y(n1396)
         );
  INVX1 U446 ( .A(n530), .Y(n172) );
  AOI2BB2X1 U447 ( .B0(n46), .B1(n433), .A0N(n1519), .A1N(n113), .Y(n1402) );
  OAI21XL U448 ( .A0(n1404), .A1(n1405), .B0(n149), .Y(n1403) );
  OAI211X1 U449 ( .A0(n122), .A1(n305), .B0(n319), .C0(n219), .Y(n317) );
  INVX1 U450 ( .A(n1366), .Y(n209) );
  AOI211X1 U451 ( .A0(n120), .A1(n146), .B0(n1317), .C0(n1325), .Y(n1366) );
  INVX1 U452 ( .A(n1113), .Y(n1435) );
  OAI211X1 U453 ( .A0(n1449), .A1(n33), .B0(n1044), .C0(n1105), .Y(n1113) );
  INVX1 U454 ( .A(n545), .Y(n189) );
  OAI211X1 U455 ( .A0(n1524), .A1(n46), .B0(n501), .C0(n537), .Y(n545) );
  INVX1 U456 ( .A(n792), .Y(n1486) );
  OAI211X1 U457 ( .A0(n1500), .A1(n59), .B0(n748), .C0(n784), .Y(n792) );
  OAI22XL U458 ( .A0(n204), .A1(n147), .B0(n190), .B1(n223), .Y(n1316) );
  NOR4X1 U459 ( .A(n1047), .B(n1048), .C(n925), .D(n1049), .Y(n1040) );
  OAI22XL U460 ( .A0(n24), .A1(n1438), .B0(n1423), .B1(n1452), .Y(n1047) );
  NOR4X1 U461 ( .A(n751), .B(n752), .C(n598), .D(n753), .Y(n744) );
  OAI22XL U462 ( .A0(n50), .A1(n1489), .B0(n1474), .B1(n1503), .Y(n751) );
  OAI21XL U463 ( .A0(n261), .A1(n1545), .B0(n262), .Y(n258) );
  NOR3X1 U464 ( .A(n1103), .B(n1100), .C(n1104), .Y(n1091) );
  OAI22XL U465 ( .A0(n43), .A1(n29), .B0(n30), .B1(n35), .Y(n1104) );
  NAND4BX1 U466 ( .AN(n1037), .B(n1105), .C(n1433), .D(n1427), .Y(n1103) );
  NOR3X1 U467 ( .A(n535), .B(n532), .C(n536), .Y(n523) );
  OAI22XL U468 ( .A0(n80), .A1(n12), .B0(n13), .B1(n72), .Y(n536) );
  NAND4BX1 U469 ( .AN(n494), .B(n537), .C(n187), .D(n181), .Y(n535) );
  NOR3X1 U470 ( .A(n782), .B(n779), .C(n783), .Y(n770) );
  OAI22XL U471 ( .A0(n69), .A1(n55), .B0(n56), .B1(n61), .Y(n783) );
  NAND4BX1 U472 ( .AN(n741), .B(n784), .C(n1484), .D(n1478), .Y(n782) );
  OAI22XL U473 ( .A0(n274), .A1(n226), .B0(n147), .B1(n223), .Y(n326) );
  OAI22XL U474 ( .A0(n135), .A1(n1506), .B0(n49), .B1(n1503), .Y(n872) );
  OAI22XL U475 ( .A0(n125), .A1(n1455), .B0(n23), .B1(n1452), .Y(n1193) );
  OAI22XL U476 ( .A0(n108), .A1(n1534), .B0(n6), .B1(n1531), .Y(n1410) );
  NAND2X1 U477 ( .A(n249), .B(n1220), .Y(n265) );
  OAI22XL U478 ( .A0(n190), .A1(n226), .B0(n222), .B1(n228), .Y(n1305) );
  OAI22XL U479 ( .A0(n1447), .A1(n23), .B0(n31), .B1(n41), .Y(n991) );
  OAI22XL U480 ( .A0(n1522), .A1(n6), .B0(n14), .B1(n78), .Y(n448) );
  OAI22XL U481 ( .A0(n1498), .A1(n49), .B0(n57), .B1(n67), .Y(n695) );
  OAI22XL U482 ( .A0(n137), .A1(n63), .B0(n1502), .B1(n52), .Y(n878) );
  OAI22XL U483 ( .A0(n127), .A1(n37), .B0(n1451), .B1(n26), .Y(n1199) );
  OAI22XL U484 ( .A0(n110), .A1(n74), .B0(n1530), .B1(n9), .Y(n1416) );
  NOR2X1 U485 ( .A(n1445), .B(n130), .Y(n1017) );
  NOR2X1 U486 ( .A(n1520), .B(n113), .Y(n474) );
  NOR2X1 U487 ( .A(n1496), .B(n140), .Y(n721) );
  NOR4BX1 U488 ( .AN(n1005), .B(n1116), .C(n1117), .D(n1046), .Y(n1107) );
  OAI222XL U489 ( .A0(n124), .A1(n1442), .B0(n1118), .B1(n28), .C0(n130), .C1(
        n1441), .Y(n1116) );
  NOR4BX1 U490 ( .AN(n462), .B(n548), .C(n549), .D(n503), .Y(n539) );
  OAI222XL U491 ( .A0(n107), .A1(n1517), .B0(n550), .B1(n11), .C0(n407), .C1(
        n1516), .Y(n548) );
  NOR4BX1 U492 ( .AN(n709), .B(n795), .C(n796), .D(n750), .Y(n786) );
  OAI222XL U493 ( .A0(n134), .A1(n1493), .B0(n797), .B1(n54), .C0(n623), .C1(
        n1492), .Y(n795) );
  NOR4X1 U494 ( .A(n504), .B(n505), .C(n382), .D(n506), .Y(n497) );
  OAI22XL U495 ( .A0(n7), .A1(n1513), .B0(n177), .B1(n1531), .Y(n504) );
  NAND2X1 U496 ( .A(n1220), .B(n88), .Y(n1255) );
  NAND2X1 U497 ( .A(n269), .B(n86), .Y(n1215) );
  NOR2X1 U498 ( .A(n1442), .B(n21), .Y(n1003) );
  NOR2X1 U499 ( .A(n1517), .B(n5), .Y(n460) );
  NOR2X1 U500 ( .A(n1493), .B(n48), .Y(n707) );
  NAND2X1 U501 ( .A(n129), .B(n973), .Y(n1000) );
  NAND2X1 U502 ( .A(n347), .B(n430), .Y(n457) );
  NAND2X1 U503 ( .A(n563), .B(n646), .Y(n704) );
  AOI211X1 U504 ( .A0(n293), .A1(n1548), .B0(n1373), .C0(n1374), .Y(n1372) );
  OAI22XL U505 ( .A0(n145), .A1(n17), .B0(n212), .B1(n143), .Y(n1374) );
  NAND4BBXL U506 ( .AN(n1232), .BN(n1349), .C(n198), .D(n1253), .Y(n1373) );
  NAND4BX1 U507 ( .AN(n1336), .B(n313), .C(n1296), .D(n1337), .Y(n1326) );
  OAI21XL U508 ( .A0(n119), .A1(n267), .B0(n121), .Y(n1337) );
  OAI222XL U509 ( .A0(n18), .A1(n268), .B0(n83), .B1(n1338), .C0(n15), .C1(n89), .Y(n1336) );
  NAND2X1 U510 ( .A(n293), .B(n85), .Y(n1315) );
  NAND4X1 U511 ( .A(n963), .B(n1148), .C(n959), .D(n1165), .Y(n1154) );
  AOI222XL U512 ( .A0(n132), .A1(n24), .B0(n890), .B1(n1016), .C0(n1007), .C1(
        n130), .Y(n1165) );
  NAND4X1 U513 ( .A(n636), .B(n827), .C(n632), .D(n844), .Y(n833) );
  AOI222XL U514 ( .A0(n576), .A1(n50), .B0(n139), .B1(n720), .C0(n711), .C1(
        n140), .Y(n844) );
  NAND4X1 U515 ( .A(n420), .B(n681), .C(n416), .D(n1078), .Y(n1067) );
  AOI222XL U516 ( .A0(n115), .A1(n7), .B0(n112), .B1(n473), .C0(n464), .C1(
        n113), .Y(n1078) );
  NAND2X1 U517 ( .A(n430), .B(n13), .Y(n422) );
  NAND2X1 U518 ( .A(n973), .B(n30), .Y(n965) );
  NAND2X1 U519 ( .A(n646), .B(n56), .Y(n638) );
  NAND2X1 U520 ( .A(n293), .B(n87), .Y(n262) );
  AOI2BB2X1 U521 ( .B0(n76), .B1(n345), .A0N(n45), .A1N(n75), .Y(n361) );
  AOI2BB2X1 U522 ( .B0(n39), .B1(n888), .A0N(n32), .A1N(n38), .Y(n904) );
  AOI2BB2X1 U523 ( .B0(n65), .B1(n561), .A0N(n58), .A1N(n64), .Y(n577) );
  NAND2X1 U524 ( .A(n126), .B(n1428), .Y(n1148) );
  NAND2X1 U525 ( .A(n136), .B(n1479), .Y(n827) );
  NAND2X1 U526 ( .A(n109), .B(n182), .Y(n681) );
  OAI21XL U527 ( .A0(n145), .A1(n305), .B0(n211), .Y(n1314) );
  OAI21XL U528 ( .A0(n415), .A1(n4), .B0(n416), .Y(n413) );
  OAI21XL U529 ( .A0(n958), .A1(n22), .B0(n959), .Y(n956) );
  OAI21XL U530 ( .A0(n631), .A1(n47), .B0(n632), .Y(n629) );
  NOR2X1 U531 ( .A(n25), .B(n1451), .Y(n1117) );
  NOR2X1 U532 ( .A(n51), .B(n1502), .Y(n796) );
  NOR2X1 U533 ( .A(n8), .B(n1530), .Y(n549) );
  BUFX2 U534 ( .A(n397), .Y(n110) );
  BUFX2 U535 ( .A(n940), .Y(n127) );
  BUFX2 U536 ( .A(n613), .Y(n137) );
  INVX1 U537 ( .A(n591), .Y(n1495) );
  INVX1 U538 ( .A(n918), .Y(n1444) );
  INVX1 U539 ( .A(n375), .Y(n1519) );
  INVX1 U540 ( .A(n1219), .Y(n194) );
  INVX1 U541 ( .A(n909), .Y(n42) );
  INVX1 U542 ( .A(n582), .Y(n68) );
  INVX1 U543 ( .A(n366), .Y(n79) );
  NOR2X1 U544 ( .A(n119), .B(n259), .Y(n1354) );
  NOR2X1 U545 ( .A(n126), .B(n131), .Y(n1118) );
  NOR2X1 U546 ( .A(n109), .B(n114), .Y(n550) );
  NOR2X1 U547 ( .A(n136), .B(n141), .Y(n797) );
  NOR2X1 U548 ( .A(n976), .B(n126), .Y(n891) );
  NOR2X1 U549 ( .A(n649), .B(n136), .Y(n564) );
  NOR2X1 U550 ( .A(n433), .B(n109), .Y(n348) );
  AND3X2 U551 ( .A(n310), .B(n1217), .C(n319), .Y(n1216) );
  NOR2X1 U552 ( .A(n191), .B(n85), .Y(n1301) );
  INVX1 U553 ( .A(n325), .Y(n214) );
  INVX1 U554 ( .A(n909), .Y(n43) );
  INVX1 U555 ( .A(n582), .Y(n69) );
  INVX1 U556 ( .A(n366), .Y(n80) );
  BUFX2 U557 ( .A(n1545), .Y(n87) );
  INVX1 U558 ( .A(n1248), .Y(n20) );
  INVX1 U559 ( .A(n328), .Y(n223) );
  INVX1 U560 ( .A(n273), .Y(n228) );
  BUFX2 U561 ( .A(n249), .Y(n116) );
  BUFX2 U562 ( .A(n267), .Y(n120) );
  NAND2X1 U563 ( .A(n44), .B(n1448), .Y(n941) );
  NAND2X1 U564 ( .A(n70), .B(n1499), .Y(n614) );
  NAND2X1 U565 ( .A(n81), .B(n1523), .Y(n398) );
  INVX1 U566 ( .A(n902), .Y(n1452) );
  INVX1 U567 ( .A(n575), .Y(n1503) );
  INVX1 U568 ( .A(n359), .Y(n1531) );
  INVX1 U569 ( .A(n2), .Y(n108) );
  INVX1 U570 ( .A(n3), .Y(n125) );
  INVX1 U571 ( .A(n1), .Y(n135) );
  INVX1 U572 ( .A(n886), .Y(n1436) );
  INVX1 U573 ( .A(n559), .Y(n1487) );
  INVX1 U574 ( .A(n343), .Y(n1456) );
  INVX1 U575 ( .A(n3), .Y(n124) );
  INVX1 U576 ( .A(n1), .Y(n134) );
  INVX1 U577 ( .A(n2), .Y(n107) );
  BUFX2 U578 ( .A(n903), .Y(n132) );
  BUFX2 U579 ( .A(n360), .Y(n115) );
  AOI211X1 U580 ( .A0(n132), .A1(n27), .B0(n1012), .C0(n1013), .Y(n1011) );
  OAI22XL U581 ( .A0(n1425), .A1(n35), .B0(n128), .B1(n1437), .Y(n1013) );
  NAND4X1 U582 ( .A(n1000), .B(n1433), .C(n896), .D(n1417), .Y(n1012) );
  AOI211X1 U583 ( .A0(n115), .A1(n10), .B0(n469), .C0(n470), .Y(n468) );
  OAI22XL U584 ( .A0(n179), .A1(n72), .B0(n111), .B1(n1512), .Y(n470) );
  NAND4X1 U585 ( .A(n457), .B(n187), .C(n353), .D(n171), .Y(n469) );
  AOI211X1 U586 ( .A0(n576), .A1(n53), .B0(n716), .C0(n717), .Y(n715) );
  OAI22XL U587 ( .A0(n1476), .A1(n61), .B0(n138), .B1(n1488), .Y(n717) );
  NAND4X1 U588 ( .A(n704), .B(n1484), .C(n569), .D(n1468), .Y(n716) );
  AOI211X1 U589 ( .A0(n107), .A1(n115), .B0(n661), .C0(n662), .Y(n657) );
  OAI22XL U590 ( .A0(n110), .A1(n1513), .B0(n345), .B1(n1514), .Y(n662) );
  OAI211X1 U591 ( .A0(n4), .A1(n1524), .B0(n462), .C0(n351), .Y(n661) );
  AOI211X1 U592 ( .A0(n124), .A1(n132), .B0(n1128), .C0(n1129), .Y(n1124) );
  OAI22XL U593 ( .A0(n127), .A1(n1438), .B0(n888), .B1(n1439), .Y(n1129) );
  OAI211X1 U594 ( .A0(n22), .A1(n1449), .B0(n1005), .C0(n894), .Y(n1128) );
  AOI211X1 U595 ( .A0(n134), .A1(n576), .B0(n807), .C0(n808), .Y(n803) );
  OAI22XL U596 ( .A0(n137), .A1(n1489), .B0(n561), .B1(n1490), .Y(n808) );
  OAI211X1 U597 ( .A0(n47), .A1(n1500), .B0(n709), .C0(n567), .Y(n807) );
  AOI211X1 U598 ( .A0(n109), .A1(n46), .B0(n659), .C0(n660), .Y(n658) );
  OAI22XL U599 ( .A0(n1520), .A1(n11), .B0(n111), .B1(n72), .Y(n660) );
  NAND4BX1 U600 ( .AN(n381), .B(n537), .C(n180), .D(n184), .Y(n659) );
  AOI211X1 U601 ( .A0(n126), .A1(n33), .B0(n1126), .C0(n1127), .Y(n1125) );
  OAI22XL U602 ( .A0(n1445), .A1(n28), .B0(n128), .B1(n35), .Y(n1127) );
  NAND4BX1 U603 ( .AN(n924), .B(n1105), .C(n1426), .D(n1430), .Y(n1126) );
  AOI211X1 U604 ( .A0(n136), .A1(n59), .B0(n805), .C0(n806), .Y(n804) );
  OAI22XL U605 ( .A0(n1496), .A1(n54), .B0(n138), .B1(n61), .Y(n806) );
  NAND4BX1 U606 ( .AN(n597), .B(n784), .C(n1477), .D(n1481), .Y(n805) );
  OAI211X1 U607 ( .A0(n309), .A1(n226), .B0(n310), .C0(n311), .Y(n301) );
  OA21XL U608 ( .A0(n312), .A1(n143), .B0(n313), .Y(n311) );
  NAND2X1 U609 ( .A(n1446), .B(n1437), .Y(n1002) );
  NAND2X1 U610 ( .A(n1497), .B(n1488), .Y(n706) );
  NAND2X1 U611 ( .A(n1521), .B(n1512), .Y(n459) );
  NAND2X1 U612 ( .A(n219), .B(n192), .Y(n308) );
  AOI211X1 U613 ( .A0(n294), .A1(n1544), .B0(n1352), .C0(n1353), .Y(n1342) );
  OAI22XL U614 ( .A0(n145), .A1(n212), .B0(n121), .B1(n191), .Y(n1353) );
  OAI211X1 U615 ( .A0(n1354), .A1(n144), .B0(n256), .C0(n1253), .Y(n1352) );
  OAI211X1 U616 ( .A0(n347), .A1(n348), .B0(n349), .C0(n350), .Y(n340) );
  AND3X2 U617 ( .A(n351), .B(n352), .C(n353), .Y(n350) );
  OAI211X1 U618 ( .A0(n129), .A1(n891), .B0(n892), .C0(n893), .Y(n883) );
  AND3X2 U619 ( .A(n894), .B(n895), .C(n896), .Y(n893) );
  OAI211X1 U620 ( .A0(n563), .A1(n564), .B0(n565), .C0(n566), .Y(n556) );
  AND3X2 U621 ( .A(n567), .B(n568), .C(n569), .Y(n566) );
  OAI211X1 U622 ( .A0(n577), .A1(n1506), .B0(n565), .C0(n863), .Y(n859) );
  AOI2BB1X1 U623 ( .A0N(n631), .A1N(n55), .B0(n765), .Y(n863) );
  OAI211X1 U624 ( .A0(n904), .A1(n1455), .B0(n892), .C0(n1184), .Y(n1180) );
  AOI2BB1X1 U625 ( .A0N(n958), .A1N(n29), .B0(n1061), .Y(n1184) );
  OAI211X1 U626 ( .A0(n361), .A1(n1534), .B0(n349), .C0(n1401), .Y(n1397) );
  AOI2BB1X1 U627 ( .A0N(n415), .A1N(n12), .B0(n518), .Y(n1401) );
  OAI211X1 U628 ( .A0(n201), .A1(n84), .B0(n335), .C0(n218), .Y(n1303) );
  OAI211X1 U629 ( .A0(n263), .A1(n1290), .B0(n335), .C0(n313), .Y(n1355) );
  AOI211X1 U630 ( .A0(n150), .A1(n370), .B0(n371), .C0(n367), .Y(n369) );
  OAI22XL U631 ( .A0(n1456), .A1(n1530), .B0(n149), .B1(n372), .Y(n371) );
  OAI211X1 U632 ( .A0(n14), .A1(n1533), .B0(n377), .C0(n174), .Y(n370) );
  NOR4X1 U633 ( .A(n373), .B(n374), .C(n375), .D(n376), .Y(n372) );
  AOI211X1 U634 ( .A0(n160), .A1(n913), .B0(n914), .C0(n910), .Y(n912) );
  OAI22XL U635 ( .A0(n1436), .A1(n1451), .B0(n159), .B1(n915), .Y(n914) );
  OAI211X1 U636 ( .A0(n31), .A1(n1454), .B0(n920), .C0(n1420), .Y(n913) );
  NOR4X1 U637 ( .A(n916), .B(n917), .C(n918), .D(n919), .Y(n915) );
  AOI211X1 U638 ( .A0(n165), .A1(n586), .B0(n587), .C0(n583), .Y(n585) );
  OAI22XL U639 ( .A0(n1487), .A1(n1502), .B0(n164), .B1(n588), .Y(n587) );
  OAI211X1 U640 ( .A0(n57), .A1(n1505), .B0(n593), .C0(n1471), .Y(n586) );
  NOR4X1 U641 ( .A(n589), .B(n590), .C(n591), .D(n592), .Y(n588) );
  INVX1 U642 ( .A(n248), .Y(n202) );
  INVX1 U643 ( .A(n240), .Y(n231) );
  INVX1 U644 ( .A(n983), .Y(n1461) );
  INVX1 U645 ( .A(n440), .Y(n1539) );
  INVX1 U646 ( .A(n687), .Y(n1511) );
  INVX1 U647 ( .A(n1302), .Y(n232) );
  OAI22XL U648 ( .A0(n92), .A1(n1514), .B0(n71), .B1(n12), .Y(n683) );
  OAI22XL U649 ( .A0(n100), .A1(n1439), .B0(n34), .B1(n29), .Y(n1150) );
  OAI22XL U650 ( .A0(n104), .A1(n1490), .B0(n60), .B1(n55), .Y(n829) );
  OAI22XL U651 ( .A0(n1547), .A1(n17), .B0(n96), .B1(n201), .Y(n1392) );
  OAI22XL U652 ( .A0(n838), .A1(n1510), .B0(n839), .B1(n1509), .Y(n834) );
  AOI211X1 U653 ( .A0(n600), .A1(n48), .B0(n840), .C0(n841), .Y(n839) );
  NOR4X1 U654 ( .A(n842), .B(n843), .C(n141), .D(n729), .Y(n838) );
  OAI222XL U655 ( .A0(n103), .A1(n1497), .B0(n50), .B1(n1503), .C0(n1505), 
        .C1(n47), .Y(n840) );
  OAI22XL U656 ( .A0(n1072), .A1(n1538), .B0(n1073), .B1(n1537), .Y(n1068) );
  AOI211X1 U657 ( .A0(n384), .A1(n5), .B0(n1074), .C0(n1075), .Y(n1073) );
  NOR4X1 U658 ( .A(n1076), .B(n1077), .C(n114), .D(n482), .Y(n1072) );
  OAI222XL U659 ( .A0(n91), .A1(n1521), .B0(n7), .B1(n1531), .C0(n1533), .C1(
        n4), .Y(n1074) );
  NOR4BX1 U660 ( .AN(n292), .B(n1260), .C(n1261), .D(n1220), .Y(n1259) );
  OAI22XL U661 ( .A0(n89), .A1(n223), .B0(n1547), .B1(n194), .Y(n1261) );
  OAI222XL U662 ( .A0(n263), .A1(n207), .B0(n95), .B1(n212), .C0(n116), .C1(
        n203), .Y(n1260) );
  NOR2X1 U663 ( .A(n224), .B(n227), .Y(n328) );
  OAI222XL U664 ( .A0(n670), .A1(n1538), .B0(n671), .B1(n1537), .C0(n672), 
        .C1(n1541), .Y(n669) );
  NOR3X1 U665 ( .A(n679), .B(n346), .C(n680), .Y(n671) );
  NOR4X1 U666 ( .A(n673), .B(n674), .C(n482), .D(n376), .Y(n672) );
  NOR4X1 U667 ( .A(n682), .B(n683), .C(n506), .D(n495), .Y(n670) );
  OAI222XL U668 ( .A0(n1137), .A1(n1460), .B0(n1138), .B1(n1459), .C0(n1139), 
        .C1(n1463), .Y(n1136) );
  NOR3X1 U669 ( .A(n1146), .B(n889), .C(n1147), .Y(n1138) );
  NOR4X1 U670 ( .A(n1140), .B(n1141), .C(n1025), .D(n919), .Y(n1139) );
  NOR4X1 U671 ( .A(n1149), .B(n1150), .C(n1049), .D(n1038), .Y(n1137) );
  OAI222XL U672 ( .A0(n1382), .A1(n230), .B0(n1383), .B1(n229), .C0(n1384), 
        .C1(n233), .Y(n1381) );
  NOR4BX1 U673 ( .AN(n1391), .B(n1392), .C(n1318), .D(n1325), .Y(n1382) );
  NOR3X1 U674 ( .A(n1390), .B(n321), .C(n1213), .Y(n1383) );
  NOR4X1 U675 ( .A(n1385), .B(n1386), .C(n260), .D(n1368), .Y(n1384) );
  OAI222XL U676 ( .A0(n816), .A1(n1510), .B0(n817), .B1(n1509), .C0(n818), 
        .C1(n1527), .Y(n815) );
  NOR3X1 U677 ( .A(n825), .B(n562), .C(n826), .Y(n817) );
  NOR4X1 U678 ( .A(n819), .B(n820), .C(n729), .D(n592), .Y(n818) );
  NOR4X1 U679 ( .A(n828), .B(n829), .C(n753), .D(n742), .Y(n816) );
  OAI22XL U680 ( .A0(n1243), .A1(n157), .B0(n154), .B1(n1244), .Y(n1239) );
  AOI211X1 U681 ( .A0(n1248), .A1(n89), .B0(n1249), .C0(n1250), .Y(n1243) );
  AOI211X1 U682 ( .A0(n289), .A1(n1245), .B0(n1246), .C0(n1247), .Y(n1244) );
  OAI22XL U683 ( .A0(n1251), .A1(n86), .B0(n312), .B1(n84), .Y(n1250) );
  OAI22XL U684 ( .A0(n1159), .A1(n1460), .B0(n1160), .B1(n1459), .Y(n1155) );
  AOI211X1 U685 ( .A0(n927), .A1(n1421), .B0(n1161), .C0(n1162), .Y(n1160) );
  NOR4X1 U686 ( .A(n1163), .B(n1164), .C(n131), .D(n1025), .Y(n1159) );
  OAI222XL U687 ( .A0(n99), .A1(n1446), .B0(n24), .B1(n1452), .C0(n1454), .C1(
        n22), .Y(n1161) );
  OAI22XL U688 ( .A0(n250), .A1(n230), .B0(n251), .B1(n229), .Y(n242) );
  AOI211X1 U689 ( .A0(n252), .A1(n85), .B0(n253), .C0(n254), .Y(n251) );
  NOR4X1 U690 ( .A(n257), .B(n258), .C(n259), .D(n260), .Y(n250) );
  OAI222XL U691 ( .A0(n94), .A1(n219), .B0(n147), .B1(n223), .C0(n225), .C1(
        n84), .Y(n253) );
  AOI211X1 U692 ( .A0(n95), .A1(n276), .B0(n1268), .C0(n328), .Y(n1389) );
  NAND2X1 U693 ( .A(n1210), .B(n95), .Y(n264) );
  INVX1 U694 ( .A(n263), .Y(n148) );
  NOR2X1 U695 ( .A(n86), .B(n95), .Y(n263) );
  NOR2X1 U696 ( .A(n117), .B(n1210), .Y(n305) );
  NOR2X1 U697 ( .A(n131), .B(n901), .Y(n887) );
  NOR2X1 U698 ( .A(n141), .B(n574), .Y(n560) );
  NOR2X1 U699 ( .A(n114), .B(n358), .Y(n344) );
  NAND2X1 U700 ( .A(n358), .B(n92), .Y(n420) );
  NAND2X1 U701 ( .A(n901), .B(n100), .Y(n963) );
  NAND2X1 U702 ( .A(n574), .B(n104), .Y(n636) );
  OAI2BB2XL U703 ( .B0(sword[15]), .B1(n1339), .A0N(sword[15]), .A1N(n1340), 
        .Y(new_sword[11]) );
  OAI222XL U704 ( .A0(n1341), .A1(n230), .B0(n1342), .B1(n229), .C0(n1343), 
        .C1(n233), .Y(n1340) );
  AOI222XL U705 ( .A0(n1356), .A1(n233), .B0(n240), .B1(n1357), .C0(n246), 
        .C1(n1358), .Y(n1339) );
  AOI221XL U706 ( .A0(n119), .A1(n249), .B0(n267), .B1(n94), .C0(n1355), .Y(
        n1341) );
  NOR2X1 U707 ( .A(n1457), .B(n1447), .Y(n903) );
  NOR2X1 U708 ( .A(n1507), .B(n1498), .Y(n576) );
  NOR2X1 U709 ( .A(n1535), .B(n1522), .Y(n360) );
  NOR2X1 U710 ( .A(n212), .B(n94), .Y(n1317) );
  NOR2X1 U711 ( .A(n1445), .B(n98), .Y(n1048) );
  NOR2X1 U712 ( .A(n1520), .B(n90), .Y(n505) );
  NOR2X1 U713 ( .A(n1496), .B(n102), .Y(n752) );
  OAI21XL U714 ( .A0(n1307), .A1(n363), .B0(n1308), .Y(new_sword[12]) );
  AOI211X1 U715 ( .A0(n246), .A1(n1326), .B0(n1327), .C0(n1328), .Y(n1307) );
  AOI22X1 U716 ( .A0(n1274), .A1(n1309), .B0(n1302), .B1(n1310), .Y(n1308) );
  AOI21X1 U717 ( .A0(n1329), .A1(n1330), .B0(n231), .Y(n1328) );
  NOR2X1 U718 ( .A(n205), .B(n225), .Y(n259) );
  NOR2X1 U719 ( .A(n96), .B(n94), .Y(n249) );
  NOR2X1 U720 ( .A(n27), .B(n101), .Y(n888) );
  NOR2X1 U721 ( .A(n10), .B(n93), .Y(n345) );
  NOR2X1 U722 ( .A(n89), .B(n94), .Y(n274) );
  NOR2X1 U723 ( .A(n53), .B(n105), .Y(n561) );
  NOR2X1 U724 ( .A(n1516), .B(n1535), .Y(n430) );
  NOR2X1 U725 ( .A(n1441), .B(n1457), .Y(n973) );
  NOR2X1 U726 ( .A(n1492), .B(n1507), .Y(n646) );
  OAI222XL U727 ( .A0(n82), .A1(n207), .B0(n116), .B1(n18), .C0(n94), .C1(n225), .Y(n1323) );
  AOI31X1 U728 ( .A0(n187), .A1(n417), .A2(n420), .B0(n151), .Y(n674) );
  AOI31X1 U729 ( .A0(n1433), .A1(n960), .A2(n963), .B0(n161), .Y(n1141) );
  AOI31X1 U730 ( .A0(n1252), .A1(n210), .A2(n264), .B0(n156), .Y(n1386) );
  AOI31X1 U731 ( .A0(n1484), .A1(n633), .A2(n636), .B0(n166), .Y(n820) );
  NAND4X1 U732 ( .A(n313), .B(n204), .C(n206), .D(n1361), .Y(n1357) );
  AOI222XL U733 ( .A0(n289), .A1(n86), .B0(n1362), .B1(n82), .C0(n249), .C1(
        n202), .Y(n1361) );
  NAND2X1 U734 ( .A(n194), .B(n192), .Y(n1362) );
  NAND4X1 U735 ( .A(n1296), .B(n207), .C(n265), .D(n1306), .Y(n1304) );
  AOI222XL U736 ( .A0(n1210), .A1(n83), .B0(n255), .B1(n89), .C0(n146), .C1(
        n276), .Y(n1306) );
  OAI221XL U737 ( .A0(n94), .A1(n1299), .B0(n15), .B1(n147), .C0(n217), .Y(
        n1297) );
  AO22X1 U738 ( .A0(n1200), .A1(n363), .B0(sword[15]), .B1(n1201), .Y(
        new_sword[15]) );
  OAI222XL U739 ( .A0(n1221), .A1(n230), .B0(n1222), .B1(n229), .C0(n1223), 
        .C1(n233), .Y(n1200) );
  OAI21XL U740 ( .A0(n1202), .A1(n233), .B0(n1203), .Y(n1201) );
  AOI221XL U741 ( .A0(n255), .A1(n118), .B0(n252), .B1(n274), .C0(n1233), .Y(
        n1221) );
  NAND2X1 U742 ( .A(n967), .B(n99), .Y(n1044) );
  NAND2X1 U743 ( .A(n424), .B(n91), .Y(n501) );
  NAND2X1 U744 ( .A(n640), .B(n103), .Y(n748) );
  NOR2X1 U745 ( .A(n967), .B(n901), .Y(n999) );
  NOR2X1 U746 ( .A(n424), .B(n358), .Y(n456) );
  NOR2X1 U747 ( .A(n640), .B(n574), .Y(n703) );
  OAI2BB2XL U748 ( .B0(n1331), .B1(n230), .A0N(n1332), .A1N(n300), .Y(n1327)
         );
  NOR4BX1 U749 ( .AN(n1315), .B(n1334), .C(n1335), .D(n260), .Y(n1331) );
  NAND4BX1 U750 ( .AN(n1333), .B(n1279), .C(n1252), .D(n292), .Y(n1332) );
  AO21X1 U751 ( .A0(n274), .A1(n1227), .B0(n1317), .Y(n1335) );
  BUFX2 U752 ( .A(n293), .Y(n119) );
  AOI211X1 U753 ( .A0(n276), .A1(n96), .B0(n1348), .C0(n1349), .Y(n1347) );
  OAI21XL U754 ( .A0(n149), .A1(n410), .B0(n411), .Y(n404) );
  AOI211X1 U755 ( .A0(n400), .A1(n396), .B0(n418), .C0(n419), .Y(n410) );
  OAI31XL U756 ( .A0(n412), .A1(n413), .A2(n414), .B0(sword[5]), .Y(n411) );
  OAI22XL U757 ( .A0(n79), .A1(n4), .B0(n182), .B1(n1514), .Y(n419) );
  OAI21XL U758 ( .A0(n159), .A1(n953), .B0(n954), .Y(n947) );
  AOI211X1 U759 ( .A0(n943), .A1(n939), .B0(n961), .C0(n962), .Y(n953) );
  OAI31XL U760 ( .A0(n955), .A1(n956), .A2(n957), .B0(sword[21]), .Y(n954) );
  OAI22XL U761 ( .A0(n42), .A1(n22), .B0(n1428), .B1(n1439), .Y(n962) );
  OAI21XL U762 ( .A0(n164), .A1(n626), .B0(n627), .Y(n620) );
  AOI211X1 U763 ( .A0(n616), .A1(n612), .B0(n634), .C0(n635), .Y(n626) );
  OAI31XL U764 ( .A0(n628), .A1(n629), .A2(n630), .B0(sword[29]), .Y(n627) );
  OAI22XL U765 ( .A0(n68), .A1(n47), .B0(n1479), .B1(n1490), .Y(n635) );
  OAI21XL U766 ( .A0(n1291), .A1(n229), .B0(n1292), .Y(n1285) );
  OAI31XL U767 ( .A0(n1293), .A1(n202), .A2(n1294), .B0(n302), .Y(n1292) );
  NOR3X1 U768 ( .A(n1297), .B(n1281), .C(n1298), .Y(n1291) );
  OAI22XL U769 ( .A0(n220), .A1(n148), .B0(n88), .B1(n207), .Y(n1294) );
  INVX1 U770 ( .A(n289), .Y(n225) );
  INVX1 U771 ( .A(n1230), .Y(n226) );
  NOR2X1 U772 ( .A(n1210), .B(n284), .Y(n1299) );
  NOR2X1 U773 ( .A(n1220), .B(n284), .Y(n1338) );
  INVX1 U774 ( .A(n378), .Y(n1534) );
  INVX1 U775 ( .A(n921), .Y(n1455) );
  INVX1 U776 ( .A(n594), .Y(n1506) );
  OAI222XL U777 ( .A0(sword[13]), .A1(n1319), .B0(n1320), .B1(n158), .C0(n228), 
        .C1(n219), .Y(n1309) );
  NOR4X1 U778 ( .A(n1321), .B(n1232), .C(n293), .D(n278), .Y(n1320) );
  NOR4X1 U779 ( .A(n1323), .B(n1324), .C(n1325), .D(n282), .Y(n1319) );
  OAI22XL U780 ( .A0(n16), .A1(n85), .B0(n190), .B1(n222), .Y(n1321) );
  BUFX2 U781 ( .A(n885), .Y(n126) );
  BUFX2 U782 ( .A(n342), .Y(n109) );
  BUFX2 U783 ( .A(n558), .Y(n136) );
  NAND2X1 U784 ( .A(n268), .B(n307), .Y(n256) );
  OAI222XL U785 ( .A0(n980), .A1(n1462), .B0(n981), .B1(n1464), .C0(n982), 
        .C1(n1465), .Y(new_sword[21]) );
  INVX1 U786 ( .A(n936), .Y(n1462) );
  AOI2BB2X1 U787 ( .B0(n1010), .B1(n162), .A0N(n1011), .A1N(n162), .Y(n981) );
  AOI221XL U788 ( .A0(n983), .A1(n984), .B0(n985), .B1(n986), .C0(n987), .Y(
        n982) );
  OAI222XL U789 ( .A0(n437), .A1(n1540), .B0(n438), .B1(n1542), .C0(n439), 
        .C1(n1543), .Y(new_sword[5]) );
  INVX1 U790 ( .A(n393), .Y(n1540) );
  AOI2BB2X1 U791 ( .B0(n467), .B1(n152), .A0N(n468), .A1N(n152), .Y(n438) );
  AOI221XL U792 ( .A0(n440), .A1(n441), .B0(n442), .B1(n443), .C0(n444), .Y(
        n439) );
  OAI222XL U793 ( .A0(n235), .A1(n236), .B0(n237), .B1(n238), .C0(sword[15]), 
        .C1(n239), .Y(new_sword[9]) );
  AOI211X1 U794 ( .A0(n240), .A1(n241), .B0(n242), .C0(n243), .Y(n239) );
  AOI222XL U795 ( .A0(n271), .A1(n157), .B0(n155), .B1(n272), .C0(n117), .C1(
        n273), .Y(n237) );
  AOI211X1 U796 ( .A0(n155), .A1(n285), .B0(n286), .C0(n287), .Y(n235) );
  OAI222XL U797 ( .A0(n684), .A1(n1526), .B0(n685), .B1(n1528), .C0(n686), 
        .C1(n1529), .Y(new_sword[29]) );
  INVX1 U798 ( .A(n609), .Y(n1526) );
  AOI2BB2X1 U799 ( .B0(n714), .B1(n167), .A0N(n715), .A1N(n167), .Y(n685) );
  AOI221XL U800 ( .A0(n687), .A1(n688), .B0(n689), .B1(n690), .C0(n691), .Y(
        n686) );
  OAI222XL U801 ( .A0(n193), .A1(sword[15]), .B0(n238), .B1(n1369), .C0(n236), 
        .C1(n1370), .Y(new_sword[10]) );
  OA22X1 U802 ( .A0(n1371), .A1(n157), .B0(n155), .B1(n1372), .Y(n1370) );
  OA22X1 U803 ( .A0(n1376), .A1(n157), .B0(n154), .B1(n1377), .Y(n1369) );
  INVX1 U804 ( .A(n1381), .Y(n193) );
  AOI211X1 U805 ( .A0(n1227), .A1(n86), .B0(n1228), .C0(n283), .Y(n1226) );
  NAND3X1 U806 ( .A(n215), .B(n194), .C(n1214), .Y(n1228) );
  NOR2X1 U807 ( .A(n1218), .B(n88), .Y(n1268) );
  INVX1 U808 ( .A(n943), .Y(n1454) );
  INVX1 U809 ( .A(n400), .Y(n1533) );
  INVX1 U810 ( .A(n616), .Y(n1505) );
  OAI22XL U811 ( .A0(n228), .A1(n191), .B0(n154), .B1(n288), .Y(n286) );
  AOI221XL U812 ( .A0(n120), .A1(n96), .B0(n274), .B1(n289), .C0(n290), .Y(
        n288) );
  OAI211X1 U813 ( .A0(n291), .A1(n82), .B0(n292), .C0(n198), .Y(n290) );
  NOR2X1 U814 ( .A(n119), .B(n294), .Y(n291) );
  INVX1 U815 ( .A(n95), .Y(n1548) );
  OAI22XL U816 ( .A0(n330), .A1(n156), .B0(n154), .B1(n331), .Y(n329) );
  AOI221XL U817 ( .A0(n307), .A1(n82), .B0(n119), .B1(n95), .C0(n334), .Y(n330) );
  AOI211X1 U818 ( .A0(n332), .A1(n144), .B0(n333), .C0(n277), .Y(n331) );
  OAI211X1 U819 ( .A0(n144), .A1(n191), .B0(n335), .C0(n18), .Y(n334) );
  INVX1 U820 ( .A(sword[2]), .Y(n75) );
  INVX1 U821 ( .A(sword[18]), .Y(n38) );
  INVX1 U822 ( .A(sword[26]), .Y(n64) );
  OAI31XL U823 ( .A0(n1204), .A1(n1205), .A2(n1206), .B0(n233), .Y(n1203) );
  OAI22XL U824 ( .A0(n309), .A1(n226), .B0(n228), .B1(n204), .Y(n1206) );
  OAI221XL U825 ( .A0(n1207), .A1(n156), .B0(n155), .B1(n1208), .C0(n292), .Y(
        n1204) );
  AOI221XL U826 ( .A0(n1210), .A1(n86), .B0(n328), .B1(sword[8]), .C0(n120), 
        .Y(n1207) );
  INVX1 U827 ( .A(n1055), .Y(n1447) );
  INVX1 U828 ( .A(n512), .Y(n1522) );
  INVX1 U829 ( .A(n759), .Y(n1498) );
  INVX1 U830 ( .A(n316), .Y(n220) );
  OAI222XL U831 ( .A0(n223), .A1(n1322), .B0(n249), .B1(n1251), .C0(n16), .C1(
        n88), .Y(n1333) );
  OAI2BB1X1 U832 ( .A0N(sword[8]), .A1N(n255), .B0(n256), .Y(n254) );
  AOI221XL U833 ( .A0(n328), .A1(n121), .B0(n1248), .B1(n147), .C0(n1378), .Y(
        n1377) );
  OAI211X1 U834 ( .A0(n118), .A1(n247), .B0(n1217), .C0(n194), .Y(n1378) );
  INVX1 U835 ( .A(n926), .Y(n1448) );
  INVX1 U836 ( .A(n383), .Y(n1523) );
  INVX1 U837 ( .A(n599), .Y(n1499) );
  INVX1 U838 ( .A(n98), .Y(n1428) );
  INVX1 U839 ( .A(n90), .Y(n182) );
  INVX1 U840 ( .A(n102), .Y(n1479) );
  INVX1 U841 ( .A(sword[8]), .Y(n1545) );
  AOI222XL U842 ( .A0(n1109), .A1(n161), .B0(n160), .B1(n1110), .C0(n886), 
        .C1(n1016), .Y(n1108) );
  NAND3BX1 U843 ( .AN(n1111), .B(n1112), .C(n1435), .Y(n1110) );
  NAND4BBXL U844 ( .AN(n1114), .BN(n1045), .C(n965), .D(n1115), .Y(n1109) );
  OAI22XL U845 ( .A0(n1447), .A1(n23), .B0(n1441), .B1(n28), .Y(n1111) );
  AOI222XL U846 ( .A0(n541), .A1(n151), .B0(n150), .B1(n542), .C0(n343), .C1(
        n473), .Y(n540) );
  NAND3BX1 U847 ( .AN(n543), .B(n544), .C(n189), .Y(n542) );
  NAND4BBXL U848 ( .AN(n546), .BN(n502), .C(n422), .D(n547), .Y(n541) );
  OAI22XL U849 ( .A0(n1522), .A1(n6), .B0(n1516), .B1(n12), .Y(n543) );
  AOI222XL U850 ( .A0(n788), .A1(n166), .B0(n165), .B1(n789), .C0(n559), .C1(
        n720), .Y(n787) );
  NAND3BX1 U851 ( .AN(n790), .B(n791), .C(n1486), .Y(n789) );
  NAND4BBXL U852 ( .AN(n793), .BN(n749), .C(n638), .D(n794), .Y(n788) );
  OAI22XL U853 ( .A0(n1498), .A1(n49), .B0(n1492), .B1(n55), .Y(n790) );
  AOI222XL U854 ( .A0(n1344), .A1(n157), .B0(n155), .B1(n1345), .C0(n269), 
        .C1(n273), .Y(n1343) );
  NAND3X1 U855 ( .A(n1346), .B(n280), .C(n1347), .Y(n1345) );
  NAND4BX1 U856 ( .AN(n1350), .B(n1315), .C(n1255), .D(n1351), .Y(n1344) );
  AOI2BB2X1 U857 ( .B0(n316), .B1(n145), .A0N(n203), .A1N(n143), .Y(n1346) );
  OAI221XL U858 ( .A0(n128), .A1(n1451), .B0(n124), .B1(n1447), .C0(n1168), 
        .Y(n1167) );
  AOI211X1 U859 ( .A0(n977), .A1(n27), .B0(n1142), .C0(n910), .Y(n1168) );
  OAI221XL U860 ( .A0(n138), .A1(n1502), .B0(n134), .B1(n1498), .C0(n847), .Y(
        n846) );
  AOI211X1 U861 ( .A0(n650), .A1(n53), .B0(n821), .C0(n583), .Y(n847) );
  OAI221XL U862 ( .A0(n111), .A1(n1530), .B0(n107), .B1(n1522), .C0(n1081), 
        .Y(n1080) );
  AOI211X1 U863 ( .A0(n434), .A1(n10), .B0(n675), .C0(n367), .Y(n1081) );
  OAI221XL U864 ( .A0(n201), .A1(n85), .B0(n225), .B1(n1546), .C0(n1267), .Y(
        n1263) );
  AOI211X1 U865 ( .A0(n307), .A1(n1245), .B0(n1242), .C0(n1268), .Y(n1267) );
  OAI221XL U866 ( .A0(n113), .A1(n1519), .B0(n110), .B1(n1531), .C0(n408), .Y(
        n406) );
  AOI211X1 U867 ( .A0(n409), .A1(n12), .B0(n382), .C0(n399), .Y(n408) );
  OAI221XL U868 ( .A0(n950), .A1(n1444), .B0(n127), .B1(n1452), .C0(n951), .Y(
        n949) );
  AOI211X1 U869 ( .A0(n952), .A1(n29), .B0(n925), .C0(n942), .Y(n951) );
  AOI222XL U870 ( .A0(n1094), .A1(n161), .B0(n160), .B1(n1095), .C0(n886), 
        .C1(n1096), .Y(n1093) );
  OAI211X1 U871 ( .A0(n891), .A1(n23), .B0(n1431), .C0(n1097), .Y(n1095) );
  NAND4BBXL U872 ( .AN(n1038), .BN(n1003), .C(n965), .D(n1099), .Y(n1094) );
  NOR2X1 U873 ( .A(n1003), .B(n1098), .Y(n1097) );
  AOI222XL U874 ( .A0(n526), .A1(n151), .B0(n150), .B1(n527), .C0(n343), .C1(
        n528), .Y(n525) );
  OAI211X1 U875 ( .A0(n348), .A1(n6), .B0(n185), .C0(n529), .Y(n527) );
  NAND4BBXL U876 ( .AN(n495), .BN(n460), .C(n422), .D(n531), .Y(n526) );
  NOR2X1 U877 ( .A(n460), .B(n530), .Y(n529) );
  AOI222XL U878 ( .A0(n773), .A1(n166), .B0(n165), .B1(n774), .C0(n559), .C1(
        n775), .Y(n772) );
  OAI211X1 U879 ( .A0(n564), .A1(n49), .B0(n1482), .C0(n776), .Y(n774) );
  NAND4BBXL U880 ( .AN(n742), .BN(n707), .C(n638), .D(n778), .Y(n773) );
  NOR2X1 U881 ( .A(n707), .B(n777), .Y(n776) );
  OAI221XL U882 ( .A0(n1269), .A1(n232), .B0(n1270), .B1(n363), .C0(n1271), 
        .Y(new_sword[13]) );
  AO21X1 U883 ( .A0(n1272), .A1(n1273), .B0(n234), .Y(n1271) );
  AOI211X1 U884 ( .A0(n246), .A1(n1284), .B0(n1285), .C0(n1286), .Y(n1270) );
  AOI221XL U885 ( .A0(n155), .A1(n1303), .B0(n1304), .B1(n156), .C0(n1305), 
        .Y(n1269) );
  AOI221XL U886 ( .A0(n581), .A1(n559), .B0(n594), .B1(n724), .C0(n725), .Y(
        n684) );
  OAI211X1 U887 ( .A0(sword[29]), .A1(n726), .B0(n727), .C0(n1470), .Y(n725)
         );
  OAI21XL U888 ( .A0(n728), .A1(n729), .B0(n164), .Y(n727) );
  INVX1 U889 ( .A(n607), .Y(n1470) );
  AOI221XL U890 ( .A0(n284), .A1(n89), .B0(n117), .B1(n143), .C0(n1209), .Y(
        n1208) );
  OAI211X1 U891 ( .A0(n118), .A1(n222), .B0(n200), .C0(n19), .Y(n1209) );
  AOI211X1 U892 ( .A0(n155), .A1(n1224), .B0(n1225), .C0(n278), .Y(n1223) );
  OAI211X1 U893 ( .A0(n225), .A1(n88), .B0(n1229), .C0(n208), .Y(n1224) );
  OAI22XL U894 ( .A0(n222), .A1(n228), .B0(n154), .B1(n1226), .Y(n1225) );
  OAI21XL U895 ( .A0(n120), .A1(n1230), .B0(n85), .Y(n1229) );
  OAI222XL U896 ( .A0(n314), .A1(n156), .B0(sword[13]), .B1(n315), .C0(n1545), 
        .C1(n219), .Y(n299) );
  AOI2BB2X1 U897 ( .B0(n89), .B1(n294), .A0N(n194), .A1N(n118), .Y(n315) );
  AOI211X1 U898 ( .A0(n268), .A1(n316), .B0(n317), .C0(n318), .Y(n314) );
  OAI22XL U899 ( .A0(n1547), .A1(n226), .B0(n274), .B1(n223), .Y(n318) );
  OAI221XL U900 ( .A0(n146), .A1(n222), .B0(n274), .B1(n220), .C0(n275), .Y(
        n272) );
  AOI211X1 U901 ( .A0(n276), .A1(n87), .B0(n277), .C0(n278), .Y(n275) );
  OAI221XL U902 ( .A0(n270), .A1(n194), .B0(n116), .B1(n223), .C0(n1241), .Y(
        n1240) );
  AOI211X1 U903 ( .A0(n255), .A1(n1547), .B0(n325), .C0(n1242), .Y(n1241) );
  OAI221XL U904 ( .A0(n140), .A1(n1495), .B0(n137), .B1(n1503), .C0(n624), .Y(
        n622) );
  AOI211X1 U905 ( .A0(n625), .A1(n55), .B0(n598), .C0(n615), .Y(n624) );
  OAI211X1 U906 ( .A0(n261), .A1(n228), .B0(n1363), .C0(n1364), .Y(n1356) );
  OAI31XL U907 ( .A0(n1367), .A1(n1301), .A2(n1368), .B0(sword[13]), .Y(n1363)
         );
  OAI21XL U908 ( .A0(n1365), .A1(n209), .B0(n157), .Y(n1364) );
  OAI21XL U909 ( .A0(n248), .A1(n87), .B0(n206), .Y(n1367) );
  AOI211X1 U910 ( .A0(n977), .A1(n128), .B0(n1026), .C0(n1027), .Y(n1022) );
  OAI211X1 U911 ( .A0(n101), .A1(n1450), .B0(n959), .C0(n41), .Y(n1026) );
  AOI211X1 U912 ( .A0(n434), .A1(n111), .B0(n483), .C0(n484), .Y(n479) );
  OAI211X1 U913 ( .A0(n93), .A1(n1525), .B0(n416), .C0(n78), .Y(n483) );
  AOI221XL U914 ( .A0(n908), .A1(n886), .B0(n921), .B1(n1020), .C0(n1021), .Y(
        n980) );
  OAI211X1 U915 ( .A0(sword[21]), .A1(n1022), .B0(n1023), .C0(n1419), .Y(n1021) );
  OAI21XL U916 ( .A0(n1024), .A1(n1025), .B0(n159), .Y(n1023) );
  INVX1 U917 ( .A(n934), .Y(n1419) );
  AOI221XL U918 ( .A0(n365), .A1(n343), .B0(n378), .B1(n477), .C0(n478), .Y(
        n437) );
  OAI211X1 U919 ( .A0(sword[5]), .A1(n479), .B0(n480), .C0(n173), .Y(n478) );
  OAI21XL U920 ( .A0(n481), .A1(n482), .B0(n149), .Y(n480) );
  INVX1 U921 ( .A(n391), .Y(n173) );
  AOI211X1 U922 ( .A0(n650), .A1(n138), .B0(n730), .C0(n731), .Y(n726) );
  OAI211X1 U923 ( .A0(n105), .A1(n1501), .B0(n632), .C0(n67), .Y(n730) );
  OAI211X1 U924 ( .A0(n228), .A1(n20), .B0(n322), .C0(n323), .Y(n320) );
  OAI31XL U925 ( .A0(n324), .A1(n117), .A2(n325), .B0(n156), .Y(n323) );
  OAI31XL U926 ( .A0(n326), .A1(n269), .A2(n327), .B0(sword[13]), .Y(n322) );
  OAI22XL U927 ( .A0(n249), .A1(n207), .B0(n268), .B1(n223), .Y(n324) );
  OAI211X1 U928 ( .A0(n68), .A1(n1487), .B0(n869), .C0(n870), .Y(n868) );
  OAI31XL U929 ( .A0(n871), .A1(n711), .A2(n598), .B0(n166), .Y(n870) );
  OAI31XL U930 ( .A0(n872), .A1(n720), .A2(n652), .B0(sword[29]), .Y(n869) );
  OAI22XL U931 ( .A0(n613), .A1(n67), .B0(n563), .B1(n1503), .Y(n871) );
  OAI211X1 U932 ( .A0(n42), .A1(n1436), .B0(n1190), .C0(n1191), .Y(n1189) );
  OAI31XL U933 ( .A0(n1192), .A1(n1007), .A2(n925), .B0(n161), .Y(n1191) );
  OAI31XL U934 ( .A0(n1193), .A1(n1016), .A2(n979), .B0(sword[21]), .Y(n1190)
         );
  OAI22XL U935 ( .A0(n940), .A1(n41), .B0(n129), .B1(n1452), .Y(n1192) );
  OAI211X1 U936 ( .A0(n79), .A1(n1456), .B0(n1407), .C0(n1408), .Y(n1406) );
  OAI31XL U937 ( .A0(n1409), .A1(n464), .A2(n382), .B0(n151), .Y(n1408) );
  OAI31XL U938 ( .A0(n1410), .A1(n473), .A2(n436), .B0(sword[5]), .Y(n1407) );
  OAI22XL U939 ( .A0(n397), .A1(n78), .B0(n347), .B1(n1531), .Y(n1409) );
  OAI22XL U940 ( .A0(n112), .A1(n78), .B0(n90), .B1(n1512), .Y(n373) );
  OAI22XL U941 ( .A0(n890), .A1(n41), .B0(n98), .B1(n1437), .Y(n916) );
  OAI22XL U942 ( .A0(n139), .A1(n67), .B0(n102), .B1(n1488), .Y(n589) );
  NOR2X1 U943 ( .A(n19), .B(sword[8]), .Y(n325) );
  NOR2X1 U944 ( .A(n205), .B(n227), .Y(n1219) );
  OAI22XL U945 ( .A0(n1056), .A1(n1460), .B0(n1057), .B1(n1459), .Y(n1051) );
  NOR4X1 U946 ( .A(n1059), .B(n1060), .C(n1025), .D(n1045), .Y(n1056) );
  NOR4BX1 U947 ( .AN(n960), .B(n1058), .C(n1017), .D(n974), .Y(n1057) );
  AO21X1 U948 ( .A0(n125), .A1(n978), .B0(n1048), .Y(n1060) );
  OAI22XL U949 ( .A0(n760), .A1(n1510), .B0(n761), .B1(n1509), .Y(n755) );
  NOR4X1 U950 ( .A(n763), .B(n764), .C(n729), .D(n749), .Y(n760) );
  NOR4BX1 U951 ( .AN(n633), .B(n762), .C(n721), .D(n647), .Y(n761) );
  AO21X1 U952 ( .A0(n135), .A1(n651), .B0(n752), .Y(n764) );
  NOR3X1 U953 ( .A(n175), .B(n152), .C(n1514), .Y(n391) );
  NOR3X1 U954 ( .A(n21), .B(n162), .C(n1439), .Y(n934) );
  NOR3X1 U955 ( .A(n1472), .B(n167), .C(n1490), .Y(n607) );
  NOR2X1 U956 ( .A(n42), .B(n99), .Y(n925) );
  NOR2X1 U957 ( .A(n68), .B(n103), .Y(n598) );
  NOR2X1 U958 ( .A(n79), .B(n91), .Y(n382) );
  OAI21XL U959 ( .A0(n98), .A1(n999), .B0(n1000), .Y(n996) );
  OAI21XL U960 ( .A0(n90), .A1(n456), .B0(n457), .Y(n453) );
  OAI21XL U961 ( .A0(n102), .A1(n703), .B0(n704), .Y(n700) );
  OAI21XL U962 ( .A0(n988), .A1(n1459), .B0(n989), .Y(n987) );
  OAI31XL U963 ( .A0(n990), .A1(n1440), .A2(n991), .B0(n945), .Y(n989) );
  NOR4X1 U964 ( .A(n995), .B(n996), .C(n997), .D(n998), .Y(n988) );
  INVX1 U965 ( .A(n992), .Y(n1440) );
  OAI21XL U966 ( .A0(n445), .A1(n1537), .B0(n446), .Y(n444) );
  OAI31XL U967 ( .A0(n447), .A1(n1515), .A2(n448), .B0(n402), .Y(n446) );
  NOR4X1 U968 ( .A(n452), .B(n453), .C(n454), .D(n455), .Y(n445) );
  INVX1 U969 ( .A(n449), .Y(n1515) );
  OAI21XL U970 ( .A0(n692), .A1(n1509), .B0(n693), .Y(n691) );
  OAI31XL U971 ( .A0(n694), .A1(n1491), .A2(n695), .B0(n618), .Y(n693) );
  NOR4X1 U972 ( .A(n699), .B(n700), .C(n701), .D(n702), .Y(n692) );
  INVX1 U973 ( .A(n696), .Y(n1491) );
  NOR2X1 U974 ( .A(n120), .B(n1210), .Y(n248) );
  NOR2X1 U975 ( .A(n162), .B(n100), .Y(n886) );
  NOR2X1 U976 ( .A(n167), .B(n104), .Y(n559) );
  NOR2X1 U977 ( .A(n152), .B(n92), .Y(n343) );
  NOR2X1 U978 ( .A(n157), .B(n96), .Y(n273) );
  NOR2X1 U979 ( .A(n1507), .B(n1504), .Y(n575) );
  NOR2X1 U980 ( .A(n1457), .B(n1453), .Y(n902) );
  NOR2X1 U981 ( .A(n1535), .B(n1532), .Y(n359) );
  NOR4X1 U982 ( .A(n428), .B(n429), .C(n430), .D(n431), .Y(n427) );
  OAI22XL U983 ( .A0(n45), .A1(n1531), .B0(n1519), .B1(n12), .Y(n429) );
  OAI222XL U984 ( .A0(n345), .A1(n78), .B0(n92), .B1(n1520), .C0(n397), .C1(
        n1516), .Y(n428) );
  NOR4X1 U985 ( .A(n971), .B(n972), .C(n973), .D(n974), .Y(n970) );
  OAI22XL U986 ( .A0(n32), .A1(n1452), .B0(n1444), .B1(n29), .Y(n972) );
  OAI222XL U987 ( .A0(n888), .A1(n41), .B0(n100), .B1(n1445), .C0(n940), .C1(
        n1441), .Y(n971) );
  NOR4X1 U988 ( .A(n644), .B(n645), .C(n646), .D(n647), .Y(n643) );
  OAI22XL U989 ( .A0(n58), .A1(n1503), .B0(n1495), .B1(n55), .Y(n645) );
  OAI222XL U990 ( .A0(n561), .A1(n67), .B0(n104), .B1(n1496), .C0(n613), .C1(
        n1492), .Y(n644) );
  NOR2X1 U991 ( .A(n132), .B(n901), .Y(n992) );
  NOR2X1 U992 ( .A(n115), .B(n358), .Y(n449) );
  NOR2X1 U993 ( .A(n142), .B(n574), .Y(n696) );
  OAI22XL U994 ( .A0(n149), .A1(n394), .B0(n395), .B1(n152), .Y(n390) );
  AOI221XL U995 ( .A0(n365), .A1(n396), .B0(n110), .B1(n398), .C0(n399), .Y(
        n395) );
  AOI221XL U996 ( .A0(n400), .A1(n12), .B0(n7), .B1(n75), .C0(n401), .Y(n394)
         );
  OAI22XL U997 ( .A0(n1534), .A1(n7), .B0(n93), .B1(n72), .Y(n401) );
  OAI22XL U998 ( .A0(n159), .A1(n937), .B0(n938), .B1(n162), .Y(n933) );
  AOI221XL U999 ( .A0(n908), .A1(n939), .B0(n127), .B1(n941), .C0(n942), .Y(
        n938) );
  AOI221XL U1000 ( .A0(n943), .A1(n29), .B0(n24), .B1(n38), .C0(n944), .Y(n937) );
  OAI22XL U1001 ( .A0(n1455), .A1(n24), .B0(n101), .B1(n35), .Y(n944) );
  OAI22XL U1002 ( .A0(n164), .A1(n610), .B0(n611), .B1(n167), .Y(n606) );
  AOI221XL U1003 ( .A0(n581), .A1(n612), .B0(n137), .B1(n614), .C0(n615), .Y(
        n611) );
  AOI221XL U1004 ( .A0(n616), .A1(n55), .B0(n50), .B1(n64), .C0(n617), .Y(n610) );
  OAI22XL U1005 ( .A0(n1506), .A1(n50), .B0(n105), .B1(n61), .Y(n617) );
  OAI22XL U1006 ( .A0(n94), .A1(n18), .B0(n145), .B1(n212), .Y(n1289) );
  OAI22XL U1007 ( .A0(n513), .A1(n1538), .B0(n514), .B1(n1537), .Y(n508) );
  NOR4X1 U1008 ( .A(n516), .B(n517), .C(n482), .D(n502), .Y(n513) );
  NOR4BX1 U1009 ( .AN(n417), .B(n515), .C(n474), .D(n431), .Y(n514) );
  AO21X1 U1010 ( .A0(n108), .A1(n435), .B0(n505), .Y(n517) );
  OAI22XL U1011 ( .A0(n93), .A1(n80), .B0(n7), .B1(n1530), .Y(n414) );
  OAI22XL U1012 ( .A0(n101), .A1(n43), .B0(n24), .B1(n1451), .Y(n957) );
  OAI22XL U1013 ( .A0(n105), .A1(n69), .B0(n50), .B1(n1502), .Y(n630) );
  OAI22XL U1014 ( .A0(n1436), .A1(n1442), .B0(n1173), .B1(n162), .Y(n1172) );
  AOI211X1 U1015 ( .A0(n125), .A1(n126), .B0(n1174), .C0(n1007), .Y(n1173) );
  OAI22XL U1016 ( .A0(n124), .A1(n1454), .B0(n890), .B1(n42), .Y(n1174) );
  OAI22XL U1017 ( .A0(n1487), .A1(n1493), .B0(n852), .B1(n167), .Y(n851) );
  AOI211X1 U1018 ( .A0(n135), .A1(n136), .B0(n853), .C0(n711), .Y(n852) );
  OAI22XL U1019 ( .A0(n134), .A1(n1505), .B0(n139), .B1(n68), .Y(n853) );
  OAI22XL U1020 ( .A0(n1456), .A1(n1517), .B0(n1086), .B1(n152), .Y(n1085) );
  AOI211X1 U1021 ( .A0(n108), .A1(n109), .B0(n1087), .C0(n464), .Y(n1086) );
  OAI22XL U1022 ( .A0(n107), .A1(n1533), .B0(n112), .B1(n79), .Y(n1087) );
  NAND2X1 U1023 ( .A(n284), .B(n84), .Y(n1279) );
  OAI222XL U1024 ( .A0(n1251), .A1(n228), .B0(n1311), .B1(n156), .C0(n155), 
        .C1(n1312), .Y(n1310) );
  AOI211X1 U1025 ( .A0(n269), .A1(n95), .B0(n1313), .C0(n1314), .Y(n1312) );
  NOR4X1 U1026 ( .A(n1316), .B(n1317), .C(n325), .D(n1318), .Y(n1311) );
  NAND4X1 U1027 ( .A(n200), .B(n1315), .C(n214), .D(n1253), .Y(n1313) );
  NOR4X1 U1028 ( .A(n1101), .B(n935), .C(n131), .D(n1061), .Y(n1092) );
  OAI221XL U1029 ( .A0(n992), .A1(n31), .B0(n99), .B1(n1454), .C0(n1102), .Y(
        n1101) );
  OAI21XL U1030 ( .A0(n978), .A1(n918), .B0(n26), .Y(n1102) );
  AOI2BB2X1 U1031 ( .B0(n205), .B1(n145), .A0N(n205), .A1N(n1548), .Y(n309) );
  NOR2X1 U1032 ( .A(n220), .B(n227), .Y(n267) );
  OAI21XL U1033 ( .A0(n1028), .A1(n1465), .B0(n1029), .Y(new_sword[20]) );
  AOI22X1 U1034 ( .A0(n936), .A1(n1030), .B0(n1009), .B1(n1031), .Y(n1029) );
  AOI211X1 U1035 ( .A0(n985), .A1(n1050), .B0(n1051), .C0(n1052), .Y(n1028) );
  OAI222XL U1036 ( .A0(n1039), .A1(n1436), .B0(n1040), .B1(n163), .C0(n160), 
        .C1(n1041), .Y(n1030) );
  OAI21XL U1037 ( .A0(n485), .A1(n1543), .B0(n486), .Y(new_sword[4]) );
  AOI22X1 U1038 ( .A0(n393), .A1(n487), .B0(n466), .B1(n488), .Y(n486) );
  AOI211X1 U1039 ( .A0(n442), .A1(n507), .B0(n508), .C0(n509), .Y(n485) );
  OAI222XL U1040 ( .A0(n496), .A1(n1456), .B0(n497), .B1(n153), .C0(n150), 
        .C1(n498), .Y(n487) );
  OAI21XL U1041 ( .A0(n732), .A1(n1529), .B0(n733), .Y(new_sword[28]) );
  AOI22X1 U1042 ( .A0(n609), .A1(n734), .B0(n713), .B1(n735), .Y(n733) );
  AOI211X1 U1043 ( .A0(n689), .A1(n754), .B0(n755), .C0(n756), .Y(n732) );
  OAI222XL U1044 ( .A0(n743), .A1(n1487), .B0(n744), .B1(n168), .C0(n165), 
        .C1(n745), .Y(n734) );
  NOR2X1 U1045 ( .A(n101), .B(n98), .Y(n940) );
  NOR2X1 U1046 ( .A(n105), .B(n102), .Y(n613) );
  NOR2X1 U1047 ( .A(n93), .B(n90), .Y(n397) );
  OAI222XL U1048 ( .A0(n41), .A1(n26), .B0(n24), .B1(n1439), .C0(n99), .C1(
        n1454), .Y(n1035) );
  OAI222XL U1049 ( .A0(n78), .A1(n9), .B0(n7), .B1(n1514), .C0(n91), .C1(n1533), .Y(n492) );
  OAI222XL U1050 ( .A0(n67), .A1(n52), .B0(n50), .B1(n1490), .C0(n103), .C1(
        n1505), .Y(n739) );
  OAI2BB1X1 U1051 ( .A0N(n1096), .A1N(n98), .B0(n1148), .Y(n1164) );
  OAI2BB1X1 U1052 ( .A0N(n775), .A1N(n102), .B0(n827), .Y(n843) );
  OAI2BB1X1 U1053 ( .A0N(n528), .A1N(n90), .B0(n681), .Y(n1077) );
  NAND2X1 U1054 ( .A(n127), .B(n909), .Y(n896) );
  NAND2X1 U1055 ( .A(n110), .B(n366), .Y(n353) );
  NAND2X1 U1056 ( .A(n137), .B(n582), .Y(n569) );
  NAND4X1 U1057 ( .A(n184), .B(n71), .C(n174), .D(n432), .Y(n426) );
  AOI222XL U1058 ( .A0(n433), .A1(n182), .B0(n434), .B1(n46), .C0(n435), .C1(
        n345), .Y(n432) );
  NAND4X1 U1059 ( .A(n1430), .B(n34), .C(n1420), .D(n975), .Y(n969) );
  AOI222XL U1060 ( .A0(n976), .A1(n1428), .B0(n977), .B1(n33), .C0(n978), .C1(
        n888), .Y(n975) );
  NAND4X1 U1061 ( .A(n1253), .B(n17), .C(n208), .D(n1262), .Y(n1258) );
  AOI222XL U1062 ( .A0(n294), .A1(n87), .B0(n276), .B1(n1548), .C0(n1227), 
        .C1(n146), .Y(n1262) );
  NAND4X1 U1063 ( .A(n1481), .B(n60), .C(n1471), .D(n648), .Y(n642) );
  AOI222XL U1064 ( .A0(n649), .A1(n1479), .B0(n650), .B1(n59), .C0(n651), .C1(
        n561), .Y(n648) );
  NOR4X1 U1065 ( .A(n533), .B(n392), .C(n114), .D(n518), .Y(n524) );
  OAI221XL U1066 ( .A0(n449), .A1(n14), .B0(n91), .B1(n1533), .C0(n534), .Y(
        n533) );
  OAI21XL U1067 ( .A0(n435), .A1(n375), .B0(n9), .Y(n534) );
  NOR4X1 U1068 ( .A(n780), .B(n608), .C(n141), .D(n765), .Y(n771) );
  OAI221XL U1069 ( .A0(n696), .A1(n57), .B0(n103), .B1(n1505), .C0(n781), .Y(
        n780) );
  OAI21XL U1070 ( .A0(n651), .A1(n591), .B0(n52), .Y(n781) );
  NAND2X1 U1071 ( .A(n1248), .B(n96), .Y(n313) );
  NAND2X1 U1072 ( .A(n424), .B(n6), .Y(n462) );
  NAND2X1 U1073 ( .A(n967), .B(n23), .Y(n1005) );
  NAND2X1 U1074 ( .A(n640), .B(n49), .Y(n709) );
  NAND4BX1 U1075 ( .AN(n421), .B(n184), .C(n422), .D(n423), .Y(n403) );
  OAI22XL U1076 ( .A0(n111), .A1(n1517), .B0(n14), .B1(n1512), .Y(n421) );
  AOI221XL U1077 ( .A0(n107), .A1(n424), .B0(n407), .B1(n378), .C0(n425), .Y(
        n423) );
  NAND4BX1 U1078 ( .AN(n964), .B(n1430), .C(n965), .D(n966), .Y(n946) );
  OAI22XL U1079 ( .A0(n128), .A1(n1442), .B0(n31), .B1(n1437), .Y(n964) );
  AOI221XL U1080 ( .A0(n124), .A1(n967), .B0(n130), .B1(n921), .C0(n968), .Y(
        n966) );
  NAND4BX1 U1081 ( .AN(n1254), .B(n1253), .C(n1255), .D(n1256), .Y(n1238) );
  OAI22XL U1082 ( .A0(n145), .A1(n191), .B0(n1546), .B1(n192), .Y(n1254) );
  AOI221XL U1083 ( .A0(n274), .A1(n284), .B0(n118), .B1(n1230), .C0(n1257), 
        .Y(n1256) );
  NAND4BX1 U1084 ( .AN(n637), .B(n1481), .C(n638), .D(n639), .Y(n619) );
  OAI22XL U1085 ( .A0(n138), .A1(n1493), .B0(n57), .B1(n1488), .Y(n637) );
  AOI221XL U1086 ( .A0(n134), .A1(n640), .B0(n623), .B1(n594), .C0(n641), .Y(
        n639) );
  NAND4BX1 U1087 ( .AN(n1061), .B(n1000), .C(n1062), .D(n1063), .Y(n1050) );
  OAI21XL U1088 ( .A0(n126), .A1(n132), .B0(n124), .Y(n1062) );
  AOI221XL U1089 ( .A0(n129), .A1(n967), .B0(n1016), .B1(n101), .C0(n1027), 
        .Y(n1063) );
  NAND4BX1 U1090 ( .AN(n518), .B(n457), .C(n519), .D(n520), .Y(n507) );
  OAI21XL U1091 ( .A0(n109), .A1(n115), .B0(n107), .Y(n519) );
  AOI221XL U1092 ( .A0(n347), .A1(n424), .B0(n473), .B1(n93), .C0(n484), .Y(
        n520) );
  NAND4BX1 U1093 ( .AN(n765), .B(n704), .C(n766), .D(n767), .Y(n754) );
  OAI21XL U1094 ( .A0(n136), .A1(n576), .B0(n134), .Y(n766) );
  AOI221XL U1095 ( .A0(n563), .A1(n640), .B0(n720), .B1(n105), .C0(n731), .Y(
        n767) );
  AOI211X1 U1096 ( .A0(n1210), .A1(n121), .B0(n1379), .C0(n1380), .Y(n1376) );
  OAI22XL U1097 ( .A0(n201), .A1(n87), .B0(n1354), .B1(n1546), .Y(n1380) );
  NAND4X1 U1098 ( .A(n1279), .B(n1215), .C(n217), .D(n215), .Y(n1379) );
  NOR2X1 U1099 ( .A(n119), .B(n1210), .Y(n1251) );
  NOR2X1 U1100 ( .A(n433), .B(n424), .Y(n415) );
  NOR2X1 U1101 ( .A(n976), .B(n967), .Y(n958) );
  NOR2X1 U1102 ( .A(n649), .B(n640), .Y(n631) );
  INVX1 U1103 ( .A(n151), .Y(n149) );
  INVX1 U1104 ( .A(n161), .Y(n159) );
  INVX1 U1105 ( .A(n166), .Y(n164) );
  NOR2X1 U1106 ( .A(n289), .B(n1219), .Y(n261) );
  NOR2X1 U1107 ( .A(n294), .B(n284), .Y(n312) );
  NAND3X1 U1108 ( .A(n848), .B(n791), .C(n849), .Y(n845) );
  AOI2BB2X1 U1109 ( .B0(n640), .B1(n139), .A0N(n1498), .A1N(n102), .Y(n848) );
  AOI211X1 U1110 ( .A0(n650), .A1(n613), .B0(n590), .C0(n741), .Y(n849) );
  OAI2BB2XL U1111 ( .B0(n164), .B1(n874), .A0N(n875), .A1N(n165), .Y(n873) );
  OAI221XL U1112 ( .A0(n1502), .A1(n139), .B0(n67), .B1(n59), .C0(n876), .Y(
        n875) );
  AOI211X1 U1113 ( .A0(n877), .A1(n54), .B0(n878), .C0(n821), .Y(n874) );
  AOI211X1 U1114 ( .A0(n135), .A1(n600), .B0(n728), .C0(n574), .Y(n876) );
  OAI2BB2XL U1115 ( .B0(n159), .B1(n1195), .A0N(n1196), .A1N(n160), .Y(n1194)
         );
  OAI221XL U1116 ( .A0(n1451), .A1(n890), .B0(n41), .B1(n33), .C0(n1197), .Y(
        n1196) );
  AOI211X1 U1117 ( .A0(n1198), .A1(n28), .B0(n1199), .C0(n1142), .Y(n1195) );
  AOI211X1 U1118 ( .A0(n125), .A1(n927), .B0(n1024), .C0(n901), .Y(n1197) );
  OAI2BB2XL U1119 ( .B0(n149), .B1(n1412), .A0N(n1413), .A1N(n150), .Y(n1411)
         );
  OAI221XL U1120 ( .A0(n1530), .A1(n112), .B0(n78), .B1(n46), .C0(n1414), .Y(
        n1413) );
  AOI211X1 U1121 ( .A0(n1415), .A1(n11), .B0(n1416), .C0(n675), .Y(n1412) );
  AOI211X1 U1122 ( .A0(n108), .A1(n384), .B0(n481), .C0(n358), .Y(n1414) );
  OAI21XL U1123 ( .A0(n115), .A1(n378), .B0(n4), .Y(n377) );
  OAI21XL U1124 ( .A0(n132), .A1(n921), .B0(n22), .Y(n920) );
  OAI21XL U1125 ( .A0(n576), .A1(n594), .B0(n47), .Y(n593) );
  INVX1 U1126 ( .A(n156), .Y(n154) );
  NAND2X1 U1127 ( .A(n145), .B(n1248), .Y(n292) );
  NOR2X1 U1128 ( .A(n126), .B(n901), .Y(n1039) );
  NOR2X1 U1129 ( .A(n109), .B(n358), .Y(n496) );
  NOR2X1 U1130 ( .A(n136), .B(n574), .Y(n743) );
  NAND2X1 U1131 ( .A(n973), .B(n101), .Y(n1105) );
  NAND2X1 U1132 ( .A(n430), .B(n93), .Y(n537) );
  NAND2X1 U1133 ( .A(n646), .B(n105), .Y(n784) );
  AOI21X1 U1134 ( .A0(n1053), .A1(n1054), .B0(n1461), .Y(n1052) );
  AOI221XL U1135 ( .A0(n967), .A1(n26), .B0(n977), .B1(n29), .C0(n1003), .Y(
        n1054) );
  AOI222XL U1136 ( .A0(n100), .A1(n1055), .B0(n973), .B1(n1428), .C0(n1007), 
        .C1(n32), .Y(n1053) );
  AOI21X1 U1137 ( .A0(n1287), .A1(n1288), .B0(n231), .Y(n1286) );
  AOI222XL U1138 ( .A0(n120), .A1(n84), .B0(n146), .B1(n259), .C0(n293), .C1(
        n96), .Y(n1287) );
  AOI211X1 U1139 ( .A0(n270), .A1(n199), .B0(n1289), .C0(n1283), .Y(n1288) );
  INVX1 U1140 ( .A(n1290), .Y(n199) );
  OAI222XL U1141 ( .A0(n121), .A1(n18), .B0(n118), .B1(n201), .C0(n95), .C1(
        n20), .Y(n1334) );
  OAI222XL U1142 ( .A0(n1452), .A1(n1020), .B0(n127), .B1(n1039), .C0(n31), 
        .C1(n1443), .Y(n1058) );
  OAI222XL U1143 ( .A0(n1531), .A1(n477), .B0(n110), .B1(n496), .C0(n14), .C1(
        n1518), .Y(n515) );
  OAI222XL U1144 ( .A0(n1503), .A1(n724), .B0(n137), .B1(n743), .C0(n57), .C1(
        n1494), .Y(n762) );
  INVX1 U1145 ( .A(n908), .Y(n1451) );
  INVX1 U1146 ( .A(n581), .Y(n1502) );
  INVX1 U1147 ( .A(n365), .Y(n1530) );
  INVX1 U1148 ( .A(n1322), .Y(n190) );
  INVX1 U1149 ( .A(n252), .Y(n191) );
  NOR2X1 U1150 ( .A(n289), .B(n1227), .Y(n247) );
  OAI222XL U1151 ( .A0(sword[21]), .A1(n1032), .B0(n1033), .B1(n163), .C0(
        n1446), .C1(n1436), .Y(n1031) );
  NOR4X1 U1152 ( .A(n1034), .B(n924), .C(n126), .D(n910), .Y(n1033) );
  NOR4X1 U1153 ( .A(n1035), .B(n1036), .C(n1037), .D(n1038), .Y(n1032) );
  OAI22XL U1154 ( .A0(n1443), .A1(n21), .B0(n1423), .B1(n1451), .Y(n1034) );
  OAI222XL U1155 ( .A0(sword[5]), .A1(n489), .B0(n490), .B1(n153), .C0(n1521), 
        .C1(n1456), .Y(n488) );
  NOR4X1 U1156 ( .A(n491), .B(n381), .C(n109), .D(n367), .Y(n490) );
  NOR4X1 U1157 ( .A(n492), .B(n493), .C(n494), .D(n495), .Y(n489) );
  OAI22XL U1158 ( .A0(n1518), .A1(n5), .B0(n177), .B1(n1530), .Y(n491) );
  OAI222XL U1159 ( .A0(sword[29]), .A1(n736), .B0(n737), .B1(n168), .C0(n1497), 
        .C1(n1487), .Y(n735) );
  NOR4X1 U1160 ( .A(n738), .B(n597), .C(n136), .D(n583), .Y(n737) );
  NOR4X1 U1161 ( .A(n739), .B(n740), .C(n741), .D(n742), .Y(n736) );
  OAI22XL U1162 ( .A0(n1494), .A1(n48), .B0(n1474), .B1(n1502), .Y(n738) );
  INVX1 U1163 ( .A(n307), .Y(n222) );
  INVX1 U1164 ( .A(n978), .Y(n1437) );
  INVX1 U1165 ( .A(n651), .Y(n1488) );
  INVX1 U1166 ( .A(n435), .Y(n1512) );
  NAND4BX1 U1167 ( .AN(n1004), .B(n896), .C(n1005), .D(n1006), .Y(n984) );
  OAI22XL U1168 ( .A0(n99), .A1(n35), .B0(n1008), .B1(n21), .Y(n1004) );
  AOI222XL U1169 ( .A0(n132), .A1(n21), .B0(n1007), .B1(n888), .C0(n126), .C1(
        n100), .Y(n1006) );
  NAND4BX1 U1170 ( .AN(n461), .B(n353), .C(n462), .D(n463), .Y(n441) );
  OAI22XL U1171 ( .A0(n91), .A1(n72), .B0(n465), .B1(n5), .Y(n461) );
  AOI222XL U1172 ( .A0(n115), .A1(n5), .B0(n464), .B1(n345), .C0(n109), .C1(
        n92), .Y(n463) );
  NAND4BX1 U1173 ( .AN(n708), .B(n569), .C(n709), .D(n710), .Y(n688) );
  OAI22XL U1174 ( .A0(n103), .A1(n61), .B0(n712), .B1(n48), .Y(n708) );
  AOI222XL U1175 ( .A0(n576), .A1(n48), .B0(n711), .B1(n561), .C0(n136), .C1(
        n104), .Y(n710) );
  INVX1 U1176 ( .A(n1020), .Y(n1423) );
  INVX1 U1177 ( .A(n477), .Y(n177) );
  INVX1 U1178 ( .A(n724), .Y(n1474) );
  NAND2X1 U1179 ( .A(n145), .B(n289), .Y(n335) );
  INVX1 U1180 ( .A(n1227), .Y(n192) );
  INVX1 U1181 ( .A(n384), .Y(n1517) );
  INVX1 U1182 ( .A(n600), .Y(n1493) );
  INVX1 U1183 ( .A(n927), .Y(n1442) );
  AOI222XL U1184 ( .A0(n1211), .A1(n157), .B0(n155), .B1(n1212), .C0(n119), 
        .C1(n273), .Y(n1202) );
  OAI221XL U1185 ( .A0(sword[8]), .A1(n305), .B0(n146), .B1(n15), .C0(n216), 
        .Y(n1212) );
  NAND4X1 U1186 ( .A(n1214), .B(n213), .C(n1215), .D(n1216), .Y(n1211) );
  INVX1 U1187 ( .A(n1213), .Y(n216) );
  AOI222XL U1188 ( .A0(n316), .A1(n96), .B0(n1220), .B1(n87), .C0(n259), .C1(
        n1548), .Y(n1329) );
  AOI21X1 U1189 ( .A0(n510), .A1(n511), .B0(n1539), .Y(n509) );
  AOI221XL U1190 ( .A0(n424), .A1(n9), .B0(n434), .B1(n12), .C0(n460), .Y(n511) );
  AOI222XL U1191 ( .A0(n92), .A1(n512), .B0(n430), .B1(n182), .C0(n464), .C1(
        n45), .Y(n510) );
  AOI21X1 U1192 ( .A0(n757), .A1(n758), .B0(n1511), .Y(n756) );
  AOI221XL U1193 ( .A0(n640), .A1(n52), .B0(n650), .B1(n55), .C0(n707), .Y(
        n758) );
  AOI222XL U1194 ( .A0(n104), .A1(n759), .B0(n646), .B1(n1479), .C0(n711), 
        .C1(n58), .Y(n757) );
  AOI221XL U1195 ( .A0(n358), .A1(n10), .B0(n359), .B1(n91), .C0(n115), .Y(
        n357) );
  AOI221XL U1196 ( .A0(n901), .A1(n27), .B0(n902), .B1(n99), .C0(n132), .Y(
        n900) );
  AOI221XL U1197 ( .A0(n574), .A1(n53), .B0(n575), .B1(n103), .C0(n576), .Y(
        n573) );
  NOR2X1 U1198 ( .A(n943), .B(n978), .Y(n1133) );
  NOR2X1 U1199 ( .A(n616), .B(n651), .Y(n812) );
  NOR2X1 U1200 ( .A(n400), .B(n435), .Y(n666) );
  AOI221XL U1201 ( .A0(n284), .A1(n83), .B0(n276), .B1(n143), .C0(n1301), .Y(
        n1330) );
  NAND3X1 U1202 ( .A(n1169), .B(n1112), .C(n1170), .Y(n1166) );
  AOI2BB2X1 U1203 ( .B0(n967), .B1(n890), .A0N(n1447), .A1N(n98), .Y(n1169) );
  AOI211X1 U1204 ( .A0(n977), .A1(n940), .B0(n917), .C0(n1037), .Y(n1170) );
  NAND3X1 U1205 ( .A(n279), .B(n280), .C(n281), .Y(n271) );
  AOI2BB2X1 U1206 ( .B0(n284), .B1(n268), .A0N(n220), .A1N(n94), .Y(n279) );
  AOI211X1 U1207 ( .A0(n116), .A1(n276), .B0(n282), .C0(n283), .Y(n281) );
  NAND3X1 U1208 ( .A(n1082), .B(n544), .C(n1083), .Y(n1079) );
  AOI2BB2X1 U1209 ( .B0(n424), .B1(n112), .A0N(n1522), .A1N(n90), .Y(n1082) );
  AOI211X1 U1210 ( .A0(n434), .A1(n397), .B0(n374), .C0(n494), .Y(n1083) );
  NAND3X1 U1211 ( .A(n861), .B(n560), .C(n862), .Y(n860) );
  AOI2BB2X1 U1212 ( .B0(n1479), .B1(n581), .A0N(n1505), .A1N(n563), .Y(n861)
         );
  AOI211X1 U1213 ( .A0(n134), .A1(n706), .B0(n701), .C0(n590), .Y(n862) );
  NAND3X1 U1214 ( .A(n1182), .B(n887), .C(n1183), .Y(n1181) );
  AOI2BB2X1 U1215 ( .B0(n1428), .B1(n908), .A0N(n1454), .A1N(n129), .Y(n1182)
         );
  AOI211X1 U1216 ( .A0(n124), .A1(n1002), .B0(n997), .C0(n917), .Y(n1183) );
  NAND3X1 U1217 ( .A(n1399), .B(n344), .C(n1400), .Y(n1398) );
  AOI2BB2X1 U1218 ( .B0(n182), .B1(n365), .A0N(n1533), .A1N(n347), .Y(n1399)
         );
  AOI211X1 U1219 ( .A0(n107), .A1(n459), .B0(n454), .C0(n374), .Y(n1400) );
  NAND3X1 U1220 ( .A(n304), .B(n305), .C(n306), .Y(n303) );
  AOI2BB2X1 U1221 ( .B0(n94), .B1(n293), .A0N(n225), .A1N(n268), .Y(n304) );
  AOI221XL U1222 ( .A0(n307), .A1(n87), .B0(n121), .B1(n308), .C0(n283), .Y(
        n306) );
  AOI211X1 U1223 ( .A0(n354), .A1(n151), .B0(n355), .C0(n356), .Y(n338) );
  OAI21XL U1224 ( .A0(n357), .A1(n151), .B0(n178), .Y(n356) );
  OAI221XL U1225 ( .A0(n1456), .A1(n1513), .B0(n361), .B1(n1534), .C0(n362), 
        .Y(n355) );
  OAI221XL U1226 ( .A0(n93), .A1(n1520), .B0(n108), .B1(n1513), .C0(n364), .Y(
        n354) );
  NAND2X1 U1227 ( .A(n599), .B(n140), .Y(n568) );
  NAND2X1 U1228 ( .A(n926), .B(n130), .Y(n895) );
  NAND2X1 U1229 ( .A(n383), .B(n113), .Y(n352) );
  AOI221XL U1230 ( .A0(n146), .A1(n1219), .B0(sword[8]), .B1(n328), .C0(n1220), 
        .Y(n310) );
  AOI211X1 U1231 ( .A0(n1016), .A1(n100), .B0(n1042), .C0(n1043), .Y(n1041) );
  OAI21XL U1232 ( .A0(n888), .A1(n887), .B0(n1044), .Y(n1043) );
  OR4X1 U1233 ( .A(n910), .B(n1045), .C(n925), .D(n1046), .Y(n1042) );
  AOI211X1 U1234 ( .A0(n473), .A1(n92), .B0(n499), .C0(n500), .Y(n498) );
  OAI21XL U1235 ( .A0(n345), .A1(n344), .B0(n501), .Y(n500) );
  OR4X1 U1236 ( .A(n367), .B(n502), .C(n382), .D(n503), .Y(n499) );
  INVX1 U1237 ( .A(sword[18]), .Y(n39) );
  INVX1 U1238 ( .A(sword[2]), .Y(n76) );
  INVX1 U1239 ( .A(sword[26]), .Y(n65) );
  NAND2X1 U1240 ( .A(n1014), .B(n1015), .Y(n1010) );
  AOI211X1 U1241 ( .A0(n977), .A1(n124), .B0(n1018), .C0(n1019), .Y(n1014) );
  NOR4X1 U1242 ( .A(n1016), .B(n925), .C(n910), .D(n1017), .Y(n1015) );
  OAI22XL U1243 ( .A0(n27), .A1(n1442), .B0(n129), .B1(n1437), .Y(n1018) );
  NAND2X1 U1244 ( .A(n471), .B(n472), .Y(n467) );
  AOI211X1 U1245 ( .A0(n434), .A1(n107), .B0(n475), .C0(n476), .Y(n471) );
  NOR4X1 U1246 ( .A(n473), .B(n382), .C(n367), .D(n474), .Y(n472) );
  OAI22XL U1247 ( .A0(n10), .A1(n1517), .B0(n347), .B1(n1512), .Y(n475) );
  NAND2X1 U1248 ( .A(n718), .B(n719), .Y(n714) );
  AOI211X1 U1249 ( .A0(n650), .A1(n134), .B0(n722), .C0(n723), .Y(n718) );
  NOR4X1 U1250 ( .A(n720), .B(n598), .C(n583), .D(n721), .Y(n719) );
  OAI22XL U1251 ( .A0(n53), .A1(n1493), .B0(n563), .B1(n1488), .Y(n722) );
  INVX1 U1252 ( .A(n300), .Y(n229) );
  INVX1 U1253 ( .A(n302), .Y(n230) );
  INVX1 U1254 ( .A(n276), .Y(n221) );
  AOI221XL U1255 ( .A0(n366), .A1(n6), .B0(n433), .B1(n9), .C0(n665), .Y(n664)
         );
  OAI221XL U1256 ( .A0(n407), .A1(n666), .B0(n1531), .B1(n11), .C0(n1519), .Y(
        n665) );
  AOI221XL U1257 ( .A0(n909), .A1(n23), .B0(n976), .B1(n26), .C0(n1132), .Y(
        n1131) );
  OAI221XL U1258 ( .A0(n130), .A1(n1133), .B0(n1452), .B1(n28), .C0(n1444), 
        .Y(n1132) );
  AOI221XL U1259 ( .A0(n582), .A1(n49), .B0(n649), .B1(n52), .C0(n811), .Y(
        n810) );
  OAI221XL U1260 ( .A0(n623), .A1(n812), .B0(n1503), .B1(n54), .C0(n1495), .Y(
        n811) );
  INVX1 U1261 ( .A(n948), .Y(n1459) );
  INVX1 U1262 ( .A(n405), .Y(n1537) );
  INVX1 U1263 ( .A(n621), .Y(n1509) );
  OR2X1 U1264 ( .A(n1218), .B(n85), .Y(n319) );
  AOI221XL U1265 ( .A0(n111), .A1(n375), .B0(n90), .B1(n359), .C0(n430), .Y(
        n349) );
  AOI221XL U1266 ( .A0(n128), .A1(n918), .B0(n98), .B1(n902), .C0(n973), .Y(
        n892) );
  AOI221XL U1267 ( .A0(n138), .A1(n591), .B0(n102), .B1(n575), .C0(n646), .Y(
        n565) );
  OAI31XL U1268 ( .A0(n1280), .A1(n1281), .A2(n1282), .B0(sword[13]), .Y(n1272) );
  OAI22XL U1269 ( .A0(sword[8]), .A1(n219), .B0(n148), .B1(n18), .Y(n1282) );
  OAI211X1 U1270 ( .A0(n263), .A1(n192), .B0(n210), .C0(n213), .Y(n1280) );
  OAI31XL U1271 ( .A0(n1275), .A1(n1276), .A2(n1277), .B0(n158), .Y(n1273) );
  OAI21XL U1272 ( .A0(n1547), .A1(n221), .B0(n1278), .Y(n1276) );
  OAI22XL U1273 ( .A0(n1545), .A1(n191), .B0(n268), .B1(n192), .Y(n1277) );
  NAND4X1 U1274 ( .A(n1279), .B(n200), .C(n214), .D(n15), .Y(n1275) );
  AOI211X1 U1275 ( .A0(n430), .A1(n90), .B0(n667), .C0(n668), .Y(n663) );
  OAI22XL U1276 ( .A0(n71), .A1(n12), .B0(n550), .B1(n14), .Y(n668) );
  NAND4BBXL U1277 ( .AN(n474), .BN(n455), .C(n351), .D(n185), .Y(n667) );
  AOI211X1 U1278 ( .A0(n973), .A1(n98), .B0(n1134), .C0(n1135), .Y(n1130) );
  OAI22XL U1279 ( .A0(n34), .A1(n29), .B0(n1118), .B1(n31), .Y(n1135) );
  NAND4BBXL U1280 ( .AN(n1017), .BN(n998), .C(n894), .D(n1431), .Y(n1134) );
  AOI211X1 U1281 ( .A0(n646), .A1(n102), .B0(n813), .C0(n814), .Y(n809) );
  OAI22XL U1282 ( .A0(n60), .A1(n55), .B0(n797), .B1(n57), .Y(n814) );
  NAND4BBXL U1283 ( .AN(n721), .BN(n702), .C(n567), .D(n1482), .Y(n813) );
  OAI221XL U1284 ( .A0(n90), .A1(n344), .B0(n345), .B1(n74), .C0(n176), .Y(
        n341) );
  INVX1 U1285 ( .A(n346), .Y(n176) );
  OAI221XL U1286 ( .A0(n98), .A1(n887), .B0(n888), .B1(n37), .C0(n1422), .Y(
        n884) );
  INVX1 U1287 ( .A(n889), .Y(n1422) );
  OAI221XL U1288 ( .A0(n102), .A1(n560), .B0(n561), .B1(n63), .C0(n1473), .Y(
        n557) );
  INVX1 U1289 ( .A(n562), .Y(n1473) );
  AOI211X1 U1290 ( .A0(n897), .A1(n161), .B0(n898), .C0(n899), .Y(n881) );
  OAI21XL U1291 ( .A0(n900), .A1(n161), .B0(n1424), .Y(n899) );
  OAI221XL U1292 ( .A0(n1436), .A1(n1438), .B0(n904), .B1(n1455), .C0(n905), 
        .Y(n898) );
  OAI221XL U1293 ( .A0(n101), .A1(n1445), .B0(n125), .B1(n1438), .C0(n907), 
        .Y(n897) );
  AOI211X1 U1294 ( .A0(n570), .A1(n166), .B0(n571), .C0(n572), .Y(n554) );
  OAI21XL U1295 ( .A0(n573), .A1(n166), .B0(n1475), .Y(n572) );
  OAI221XL U1296 ( .A0(n1487), .A1(n1489), .B0(n577), .B1(n1506), .C0(n578), 
        .Y(n571) );
  OAI221XL U1297 ( .A0(n105), .A1(n1496), .B0(n135), .B1(n1489), .C0(n580), 
        .Y(n570) );
  INVX1 U1298 ( .A(n945), .Y(n1460) );
  INVX1 U1299 ( .A(n402), .Y(n1538) );
  INVX1 U1300 ( .A(n618), .Y(n1510) );
  AO21X1 U1301 ( .A0(n99), .A1(n952), .B0(n1117), .Y(n1162) );
  AO21X1 U1302 ( .A0(n103), .A1(n625), .B0(n796), .Y(n841) );
  AO21X1 U1303 ( .A0(n91), .A1(n409), .B0(n549), .Y(n1075) );
  AOI221XL U1304 ( .A0(n345), .A1(n383), .B0(n384), .B1(n108), .C0(n385), .Y(
        n368) );
  OAI211X1 U1305 ( .A0(n5), .A1(n1525), .B0(n386), .C0(n1516), .Y(n385) );
  OAI21XL U1306 ( .A0(n365), .A1(n375), .B0(n7), .Y(n386) );
  INVX1 U1307 ( .A(n434), .Y(n1524) );
  INVX1 U1308 ( .A(n977), .Y(n1449) );
  INVX1 U1309 ( .A(n650), .Y(n1500) );
  OAI211X1 U1310 ( .A0(n940), .A1(n1448), .B0(n993), .C0(n994), .Y(n990) );
  OAI21XL U1311 ( .A0(n927), .A1(n976), .B0(n99), .Y(n993) );
  OAI211X1 U1312 ( .A0(n397), .A1(n1523), .B0(n450), .C0(n451), .Y(n447) );
  OAI21XL U1313 ( .A0(n384), .A1(n433), .B0(n91), .Y(n450) );
  OAI211X1 U1314 ( .A0(n249), .A1(n1218), .B0(n1295), .C0(n1296), .Y(n1293) );
  OAI21XL U1315 ( .A0(n252), .A1(n294), .B0(sword[8]), .Y(n1295) );
  OAI211X1 U1316 ( .A0(n613), .A1(n1499), .B0(n697), .C0(n698), .Y(n694) );
  OAI21XL U1317 ( .A0(n600), .A1(n649), .B0(n103), .Y(n697) );
  AOI211X1 U1318 ( .A0(n720), .A1(n104), .B0(n746), .C0(n747), .Y(n745) );
  OAI21XL U1319 ( .A0(n561), .A1(n560), .B0(n748), .Y(n747) );
  OR4X1 U1320 ( .A(n583), .B(n749), .C(n598), .D(n750), .Y(n746) );
  AOI211X1 U1321 ( .A0(n365), .A1(n5), .B0(n366), .C0(n367), .Y(n364) );
  AOI211X1 U1322 ( .A0(n908), .A1(n21), .B0(n909), .C0(n910), .Y(n907) );
  AOI211X1 U1323 ( .A0(n581), .A1(n48), .B0(n582), .C0(n583), .Y(n580) );
  AOI221XL U1324 ( .A0(n888), .A1(n926), .B0(n927), .B1(n125), .C0(n928), .Y(
        n911) );
  OAI211X1 U1325 ( .A0(n22), .A1(n1450), .B0(n929), .C0(n1441), .Y(n928) );
  OAI21XL U1326 ( .A0(n908), .A1(n918), .B0(n24), .Y(n929) );
  AOI221XL U1327 ( .A0(n561), .A1(n599), .B0(n600), .B1(n135), .C0(n601), .Y(
        n584) );
  OAI211X1 U1328 ( .A0(n48), .A1(n1501), .B0(n602), .C0(n1492), .Y(n601) );
  OAI21XL U1329 ( .A0(n581), .A1(n591), .B0(n50), .Y(n602) );
  OAI211X1 U1330 ( .A0(n148), .A1(n1218), .B0(n1234), .C0(n203), .Y(n1233) );
  OAI21XL U1331 ( .A0(n307), .A1(n1219), .B0(n148), .Y(n1234) );
  OAI211X1 U1332 ( .A0(n1428), .A1(n1457), .B0(n1434), .C0(n1001), .Y(n986) );
  INVX1 U1333 ( .A(n968), .Y(n1434) );
  AOI221XL U1334 ( .A0(n921), .A1(n22), .B0(n1002), .B1(n33), .C0(n1003), .Y(
        n1001) );
  OAI211X1 U1335 ( .A0(n182), .A1(n1535), .B0(n188), .C0(n458), .Y(n443) );
  INVX1 U1336 ( .A(n425), .Y(n188) );
  AOI221XL U1337 ( .A0(n378), .A1(n4), .B0(n459), .B1(n46), .C0(n460), .Y(n458) );
  OAI211X1 U1338 ( .A0(n1479), .A1(n1507), .B0(n1485), .C0(n705), .Y(n690) );
  INVX1 U1339 ( .A(n641), .Y(n1485) );
  AOI221XL U1340 ( .A0(n594), .A1(n47), .B0(n706), .B1(n59), .C0(n707), .Y(
        n705) );
  OAI211X1 U1341 ( .A0(n144), .A1(n207), .B0(n204), .C0(n295), .Y(n285) );
  AOI2BB2X1 U1342 ( .B0(n289), .B1(n143), .A0N(n20), .A1N(n268), .Y(n295) );
  OAI211X1 U1343 ( .A0(n227), .A1(n87), .B0(n197), .C0(n1300), .Y(n1284) );
  INVX1 U1344 ( .A(n1257), .Y(n197) );
  AOI221XL U1345 ( .A0(n1230), .A1(n85), .B0(n308), .B1(n89), .C0(n1301), .Y(
        n1300) );
  INVX1 U1346 ( .A(n409), .Y(n1525) );
  INVX1 U1347 ( .A(n952), .Y(n1450) );
  INVX1 U1348 ( .A(n625), .Y(n1501) );
  INVX1 U1349 ( .A(n156), .Y(n155) );
  INVX1 U1350 ( .A(n379), .Y(n169) );
  OAI221XL U1351 ( .A0(n74), .A1(n92), .B0(n1516), .B1(n347), .C0(n380), .Y(
        n379) );
  AOI211X1 U1352 ( .A0(n76), .A1(n108), .B0(n381), .C0(n382), .Y(n380) );
  INVX1 U1353 ( .A(n922), .Y(n579) );
  OAI221XL U1354 ( .A0(n37), .A1(n100), .B0(n1441), .B1(n129), .C0(n923), .Y(
        n922) );
  AOI211X1 U1355 ( .A0(n39), .A1(n125), .B0(n924), .C0(n925), .Y(n923) );
  INVX1 U1356 ( .A(n595), .Y(n1466) );
  OAI221XL U1357 ( .A0(n63), .A1(n104), .B0(n1492), .B1(n563), .C0(n596), .Y(
        n595) );
  AOI211X1 U1358 ( .A0(n65), .A1(n135), .B0(n597), .C0(n598), .Y(n596) );
  NOR2X1 U1359 ( .A(n233), .B(n97), .Y(n1302) );
  NOR2X1 U1360 ( .A(n1463), .B(n162), .Y(n985) );
  NOR2X1 U1361 ( .A(n1541), .B(n152), .Y(n442) );
  NOR2X1 U1362 ( .A(n1527), .B(n167), .Y(n689) );
  NOR2X1 U1363 ( .A(n233), .B(n154), .Y(n240) );
  NOR2X1 U1364 ( .A(n1463), .B(n159), .Y(n983) );
  NOR2X1 U1365 ( .A(n1527), .B(n164), .Y(n687) );
  NOR2X1 U1366 ( .A(n1541), .B(n149), .Y(n440) );
  NOR2X1 U1367 ( .A(n233), .B(n157), .Y(n246) );
  NAND2X1 U1368 ( .A(n97), .B(n233), .Y(n238) );
  INVX1 U1369 ( .A(n161), .Y(n160) );
  INVX1 U1370 ( .A(n166), .Y(n165) );
  INVX1 U1371 ( .A(n151), .Y(n150) );
  INVX1 U1372 ( .A(n1274), .Y(n234) );
  INVX1 U1373 ( .A(n1009), .Y(n1464) );
  INVX1 U1374 ( .A(n466), .Y(n1542) );
  INVX1 U1375 ( .A(n713), .Y(n1528) );
  INVX1 U1376 ( .A(n97), .Y(n363) );
  OAI22XL U1377 ( .A0(n228), .A1(n15), .B0(n154), .B1(n1387), .Y(n1385) );
  AOI211X1 U1378 ( .A0(sword[11]), .A1(n84), .B0(n195), .C0(n1388), .Y(n1387)
         );
  INVX1 U1379 ( .A(n1389), .Y(n195) );
  OAI22XL U1380 ( .A0(n15), .A1(n82), .B0(n95), .B1(n194), .Y(n1388) );
  OAI22XL U1381 ( .A0(n63), .A1(n1487), .B0(n164), .B1(n822), .Y(n819) );
  AOI211X1 U1382 ( .A0(sword[27]), .A1(n47), .B0(n823), .C0(n824), .Y(n822) );
  OAI221XL U1383 ( .A0(n57), .A1(n1499), .B0(n58), .B1(n1500), .C0(n1503), .Y(
        n823) );
  OAI22XL U1384 ( .A0(n1494), .A1(n52), .B0(n104), .B1(n1495), .Y(n824) );
  NOR2X1 U1385 ( .A(sword[3]), .B(sword[4]), .Y(n378) );
  NOR2X1 U1386 ( .A(sword[19]), .B(sword[20]), .Y(n921) );
  NOR2X1 U1387 ( .A(sword[27]), .B(sword[28]), .Y(n594) );
  NOR2X1 U1388 ( .A(sword[11]), .B(sword[12]), .Y(n1230) );
  NOR2X1 U1389 ( .A(sword[10]), .B(sword[12]), .Y(n276) );
  NOR2X1 U1390 ( .A(n1457), .B(sword[18]), .Y(n926) );
  NOR2X1 U1391 ( .A(n1507), .B(sword[26]), .Y(n599) );
  NOR2X1 U1392 ( .A(n1535), .B(sword[2]), .Y(n383) );
  NOR2X1 U1393 ( .A(n224), .B(sword[10]), .Y(n316) );
  NOR2X1 U1394 ( .A(n1453), .B(sword[18]), .Y(n1055) );
  NOR2X1 U1395 ( .A(n1532), .B(sword[2]), .Y(n512) );
  NOR2X1 U1396 ( .A(n1504), .B(sword[26]), .Y(n759) );
  NOR2X1 U1397 ( .A(n1455), .B(sword[18]), .Y(n885) );
  NOR2X1 U1398 ( .A(n1534), .B(sword[2]), .Y(n342) );
  NOR2X1 U1399 ( .A(n226), .B(sword[10]), .Y(n293) );
  NOR2X1 U1400 ( .A(n1506), .B(sword[26]), .Y(n558) );
  INVX1 U1401 ( .A(sword[11]), .Y(n224) );
  INVX1 U1402 ( .A(sword[27]), .Y(n1504) );
  INVX1 U1403 ( .A(sword[19]), .Y(n1453) );
  INVX1 U1404 ( .A(sword[3]), .Y(n1532) );
  BUFX2 U1405 ( .A(sword[16]), .Y(n98) );
  BUFX2 U1406 ( .A(sword[0]), .Y(n90) );
  BUFX2 U1407 ( .A(sword[24]), .Y(n102) );
  BUFX2 U1408 ( .A(sword[9]), .Y(n95) );
  BUFX2 U1409 ( .A(sword[25]), .Y(n104) );
  BUFX2 U1410 ( .A(sword[1]), .Y(n92) );
  BUFX2 U1411 ( .A(sword[17]), .Y(n100) );
  AO22X1 U1412 ( .A0(sword[23]), .A1(n1089), .B0(n1090), .B1(n1465), .Y(
        new_sword[19]) );
  OAI222XL U1413 ( .A0(n1091), .A1(n1458), .B0(n1092), .B1(n1461), .C0(
        sword[22]), .C1(n1093), .Y(n1090) );
  OAI222XL U1414 ( .A0(n1106), .A1(n1460), .B0(n1107), .B1(n1459), .C0(n1108), 
        .C1(n1463), .Y(n1089) );
  INVX1 U1415 ( .A(n985), .Y(n1458) );
  AO22X1 U1416 ( .A0(sword[7]), .A1(n521), .B0(n522), .B1(n1543), .Y(
        new_sword[3]) );
  OAI222XL U1417 ( .A0(n523), .A1(n1536), .B0(n524), .B1(n1539), .C0(sword[6]), 
        .C1(n525), .Y(n522) );
  OAI222XL U1418 ( .A0(n538), .A1(n1538), .B0(n539), .B1(n1537), .C0(n540), 
        .C1(n1541), .Y(n521) );
  INVX1 U1419 ( .A(n442), .Y(n1536) );
  AO22X1 U1420 ( .A0(sword[31]), .A1(n768), .B0(n769), .B1(n1529), .Y(
        new_sword[27]) );
  OAI222XL U1421 ( .A0(n770), .A1(n1508), .B0(n771), .B1(n1511), .C0(sword[30]), .C1(n772), .Y(n769) );
  OAI222XL U1422 ( .A0(n785), .A1(n1510), .B0(n786), .B1(n1509), .C0(n787), 
        .C1(n1527), .Y(n768) );
  INVX1 U1423 ( .A(n689), .Y(n1508) );
  BUFX2 U1424 ( .A(sword[9]), .Y(n96) );
  OAI222XL U1425 ( .A0(n296), .A1(n236), .B0(n297), .B1(n238), .C0(sword[15]), 
        .C1(n298), .Y(new_sword[8]) );
  AOI211X1 U1426 ( .A0(n269), .A1(n1548), .B0(n320), .C0(n321), .Y(n297) );
  AOI221XL U1427 ( .A0(n328), .A1(n143), .B0(n273), .B1(n284), .C0(n329), .Y(
        n296) );
  AOI222XL U1428 ( .A0(sword[14]), .A1(n299), .B0(n300), .B1(n301), .C0(n302), 
        .C1(n303), .Y(n298) );
  OAI222XL U1429 ( .A0(n1235), .A1(n232), .B0(n1236), .B1(n234), .C0(n1237), 
        .C1(n363), .Y(new_sword[14]) );
  AOI221XL U1430 ( .A0(n155), .A1(n1263), .B0(n1264), .B1(n156), .C0(n1265), 
        .Y(n1235) );
  AOI2BB2X1 U1431 ( .B0(n154), .B1(n1258), .A0N(n154), .A1N(n1259), .Y(n1236)
         );
  AOI222XL U1432 ( .A0(n302), .A1(n1238), .B0(sword[14]), .B1(n1239), .C0(n300), .C1(n1240), .Y(n1237) );
  OAI222XL U1433 ( .A0(n1151), .A1(n1122), .B0(n1152), .B1(n1120), .C0(
        sword[23]), .C1(n1153), .Y(new_sword[17]) );
  AOI211X1 U1434 ( .A0(n1171), .A1(n163), .B0(n1172), .C0(n998), .Y(n1151) );
  AOI211X1 U1435 ( .A0(n983), .A1(n1154), .B0(n1155), .C0(n1156), .Y(n1153) );
  AOI222XL U1436 ( .A0(n1166), .A1(n161), .B0(n160), .B1(n1167), .C0(n1007), 
        .C1(n886), .Y(n1152) );
  OAI222XL U1437 ( .A0(n830), .A1(n801), .B0(n831), .B1(n799), .C0(sword[31]), 
        .C1(n832), .Y(new_sword[25]) );
  AOI211X1 U1438 ( .A0(n850), .A1(n168), .B0(n851), .C0(n702), .Y(n830) );
  AOI211X1 U1439 ( .A0(n687), .A1(n833), .B0(n834), .C0(n835), .Y(n832) );
  AOI222XL U1440 ( .A0(n845), .A1(n166), .B0(n165), .B1(n846), .C0(n711), .C1(
        n559), .Y(n831) );
  OAI222XL U1441 ( .A0(n1064), .A1(n655), .B0(n1065), .B1(n653), .C0(sword[7]), 
        .C1(n1066), .Y(new_sword[1]) );
  AOI211X1 U1442 ( .A0(n1084), .A1(n153), .B0(n1085), .C0(n455), .Y(n1064) );
  AOI211X1 U1443 ( .A0(n440), .A1(n1067), .B0(n1068), .C0(n1069), .Y(n1066) );
  AOI222XL U1444 ( .A0(n1079), .A1(n151), .B0(n150), .B1(n1080), .C0(n464), 
        .C1(n343), .Y(n1065) );
  OAI222XL U1445 ( .A0(n170), .A1(sword[7]), .B0(n653), .B1(n654), .C0(n655), 
        .C1(n656), .Y(new_sword[2]) );
  OA22X1 U1446 ( .A0(n657), .A1(n152), .B0(n150), .B1(n658), .Y(n656) );
  OA22X1 U1447 ( .A0(n663), .A1(n152), .B0(n150), .B1(n664), .Y(n654) );
  INVX1 U1448 ( .A(n669), .Y(n170) );
  OAI222XL U1449 ( .A0(n906), .A1(sword[23]), .B0(n1120), .B1(n1121), .C0(
        n1122), .C1(n1123), .Y(new_sword[18]) );
  OA22X1 U1450 ( .A0(n1124), .A1(n162), .B0(n160), .B1(n1125), .Y(n1123) );
  OA22X1 U1451 ( .A0(n1130), .A1(n162), .B0(n160), .B1(n1131), .Y(n1121) );
  INVX1 U1452 ( .A(n1136), .Y(n906) );
  OAI222XL U1453 ( .A0(n1467), .A1(sword[31]), .B0(n799), .B1(n800), .C0(n801), 
        .C1(n802), .Y(new_sword[26]) );
  OA22X1 U1454 ( .A0(n803), .A1(n167), .B0(n165), .B1(n804), .Y(n802) );
  OA22X1 U1455 ( .A0(n809), .A1(n167), .B0(n165), .B1(n810), .Y(n800) );
  INVX1 U1456 ( .A(n815), .Y(n1467) );
  BUFX2 U1457 ( .A(sword[8]), .Y(n94) );
  OAI22XL U1458 ( .A0(n74), .A1(n1456), .B0(n149), .B1(n676), .Y(n673) );
  AOI211X1 U1459 ( .A0(sword[3]), .A1(n4), .B0(n677), .C0(n678), .Y(n676) );
  OAI221XL U1460 ( .A0(n14), .A1(n1523), .B0(n45), .B1(n1524), .C0(n1531), .Y(
        n677) );
  OAI22XL U1461 ( .A0(n1518), .A1(n9), .B0(n92), .B1(n1519), .Y(n678) );
  OAI22XL U1462 ( .A0(n37), .A1(n1436), .B0(n159), .B1(n1143), .Y(n1140) );
  AOI211X1 U1463 ( .A0(sword[19]), .A1(n22), .B0(n1144), .C0(n1145), .Y(n1143)
         );
  OAI221XL U1464 ( .A0(n31), .A1(n1448), .B0(n32), .B1(n1449), .C0(n1452), .Y(
        n1144) );
  OAI22XL U1465 ( .A0(n1443), .A1(n26), .B0(n100), .B1(n1444), .Y(n1145) );
  OAI221XL U1466 ( .A0(n387), .A1(n1542), .B0(n388), .B1(n1543), .C0(n389), 
        .Y(new_sword[6]) );
  OAI31XL U1467 ( .A0(n390), .A1(n391), .A2(n392), .B0(n393), .Y(n389) );
  AOI2BB2X1 U1468 ( .B0(n149), .B1(n426), .A0N(n150), .A1N(n427), .Y(n387) );
  AOI222XL U1469 ( .A0(n402), .A1(n403), .B0(sword[6]), .B1(n404), .C0(n405), 
        .C1(n406), .Y(n388) );
  OAI221XL U1470 ( .A0(n930), .A1(n1464), .B0(n931), .B1(n1465), .C0(n932), 
        .Y(new_sword[22]) );
  OAI31XL U1471 ( .A0(n933), .A1(n934), .A2(n935), .B0(n936), .Y(n932) );
  AOI2BB2X1 U1472 ( .B0(n159), .B1(n969), .A0N(n160), .A1N(n970), .Y(n930) );
  AOI222XL U1473 ( .A0(n945), .A1(n946), .B0(sword[22]), .B1(n947), .C0(n948), 
        .C1(n949), .Y(n931) );
  OAI221XL U1474 ( .A0(n603), .A1(n1528), .B0(n604), .B1(n1529), .C0(n605), 
        .Y(new_sword[30]) );
  OAI31XL U1475 ( .A0(n606), .A1(n607), .A2(n608), .B0(n609), .Y(n605) );
  AOI2BB2X1 U1476 ( .B0(n164), .B1(n642), .A0N(n165), .A1N(n643), .Y(n603) );
  AOI222XL U1477 ( .A0(n618), .A1(n619), .B0(sword[30]), .B1(n620), .C0(n621), 
        .C1(n622), .Y(n604) );
  OAI222XL U1478 ( .A0(n855), .A1(n801), .B0(n856), .B1(n799), .C0(sword[31]), 
        .C1(n857), .Y(new_sword[24]) );
  AOI221XL U1479 ( .A0(n575), .A1(n1), .B0(n640), .B1(n559), .C0(n873), .Y(
        n855) );
  AOI222XL U1480 ( .A0(sword[30]), .A1(n858), .B0(n621), .B1(n859), .C0(n618), 
        .C1(n860), .Y(n857) );
  AOI211X1 U1481 ( .A0(n720), .A1(n58), .B0(n868), .C0(n826), .Y(n856) );
  OAI222XL U1482 ( .A0(n1176), .A1(n1122), .B0(n1177), .B1(n1120), .C0(
        sword[23]), .C1(n1178), .Y(new_sword[16]) );
  AOI221XL U1483 ( .A0(n902), .A1(n28), .B0(n967), .B1(n886), .C0(n1194), .Y(
        n1176) );
  AOI222XL U1484 ( .A0(sword[22]), .A1(n1179), .B0(n948), .B1(n1180), .C0(n945), .C1(n1181), .Y(n1178) );
  AOI211X1 U1485 ( .A0(n1016), .A1(n32), .B0(n1189), .C0(n1147), .Y(n1177) );
  OAI222XL U1486 ( .A0(n1393), .A1(n655), .B0(n1394), .B1(n653), .C0(sword[7]), 
        .C1(n1395), .Y(new_sword[0]) );
  AOI221XL U1487 ( .A0(n359), .A1(n2), .B0(n424), .B1(n343), .C0(n1411), .Y(
        n1393) );
  AOI222XL U1488 ( .A0(sword[6]), .A1(n1396), .B0(n405), .B1(n1397), .C0(n402), 
        .C1(n1398), .Y(n1395) );
  AOI211X1 U1489 ( .A0(n473), .A1(n45), .B0(n1406), .C0(n680), .Y(n1394) );
  NOR2X1 U1490 ( .A(n1447), .B(sword[20]), .Y(n909) );
  NOR2X1 U1491 ( .A(n1498), .B(sword[28]), .Y(n582) );
  NOR2X1 U1492 ( .A(n1522), .B(sword[4]), .Y(n366) );
  NOR2X1 U1493 ( .A(n65), .B(sword[28]), .Y(n600) );
  NOR2X1 U1494 ( .A(n76), .B(sword[4]), .Y(n384) );
  NOR2X1 U1495 ( .A(n39), .B(sword[20]), .Y(n927) );
  NOR2X1 U1496 ( .A(n205), .B(sword[12]), .Y(n252) );
  NOR2X1 U1497 ( .A(sword[18]), .B(sword[20]), .Y(n977) );
  NOR2X1 U1498 ( .A(sword[2]), .B(sword[4]), .Y(n434) );
  NOR2X1 U1499 ( .A(sword[26]), .B(sword[28]), .Y(n650) );
  NOR2X1 U1500 ( .A(n157), .B(sword[14]), .Y(n300) );
  NOR2X1 U1501 ( .A(sword[18]), .B(sword[19]), .Y(n952) );
  NOR2X1 U1502 ( .A(sword[26]), .B(sword[27]), .Y(n625) );
  NOR2X1 U1503 ( .A(sword[2]), .B(sword[3]), .Y(n409) );
  NOR2X1 U1504 ( .A(n154), .B(sword[14]), .Y(n302) );
  NOR2X1 U1505 ( .A(n159), .B(sword[22]), .Y(n945) );
  NOR2X1 U1506 ( .A(n164), .B(sword[30]), .Y(n618) );
  NOR2X1 U1507 ( .A(n149), .B(sword[6]), .Y(n402) );
  NOR2X1 U1508 ( .A(n162), .B(sword[22]), .Y(n948) );
  NOR2X1 U1509 ( .A(n167), .B(sword[30]), .Y(n621) );
  NOR2X1 U1510 ( .A(n152), .B(sword[6]), .Y(n405) );
  NOR4BX1 U1511 ( .AN(n1217), .B(n1231), .C(n325), .D(n1232), .Y(n1222) );
  OAI22XL U1512 ( .A0(n95), .A1(n16), .B0(sword[10]), .B1(n143), .Y(n1231) );
  NAND2X1 U1513 ( .A(sword[12]), .B(n205), .Y(n1218) );
  BUFX2 U1514 ( .A(n153), .Y(n151) );
  BUFX2 U1515 ( .A(n168), .Y(n166) );
  BUFX2 U1516 ( .A(n163), .Y(n161) );
  BUFX2 U1517 ( .A(n158), .Y(n156) );
  OAI21XL U1518 ( .A0(sword[2]), .A1(n113), .B0(n11), .Y(n396) );
  OAI21XL U1519 ( .A0(sword[18]), .A1(n130), .B0(n28), .Y(n939) );
  OAI21XL U1520 ( .A0(sword[26]), .A1(n140), .B0(n54), .Y(n612) );
  BUFX2 U1521 ( .A(n163), .Y(n162) );
  BUFX2 U1522 ( .A(n153), .Y(n152) );
  BUFX2 U1523 ( .A(n168), .Y(n167) );
  OAI21XL U1524 ( .A0(sword[10]), .A1(n118), .B0(n143), .Y(n1245) );
  NOR2X1 U1525 ( .A(sword[10]), .B(sword[11]), .Y(n255) );
  BUFX2 U1526 ( .A(n158), .Y(n157) );
  BUFX2 U1527 ( .A(sword[16]), .Y(n99) );
  BUFX2 U1528 ( .A(sword[24]), .Y(n103) );
  BUFX2 U1529 ( .A(sword[0]), .Y(n91) );
  BUFX2 U1530 ( .A(sword[1]), .Y(n93) );
  BUFX2 U1531 ( .A(sword[17]), .Y(n101) );
  BUFX2 U1532 ( .A(sword[25]), .Y(n105) );
  AO22X1 U1533 ( .A0(n336), .A1(n1543), .B0(sword[7]), .B1(n337), .Y(
        new_sword[7]) );
  OAI22XL U1534 ( .A0(sword[6]), .A1(n338), .B0(n339), .B1(n1541), .Y(n337) );
  OAI222XL U1535 ( .A0(n368), .A1(n1538), .B0(n169), .B1(n1537), .C0(n369), 
        .C1(n1541), .Y(n336) );
  AOI222XL U1536 ( .A0(n340), .A1(n151), .B0(n150), .B1(n341), .C0(n109), .C1(
        n343), .Y(n339) );
  AO22X1 U1537 ( .A0(n879), .A1(n1465), .B0(sword[23]), .B1(n880), .Y(
        new_sword[23]) );
  OAI22XL U1538 ( .A0(sword[22]), .A1(n881), .B0(n882), .B1(n1463), .Y(n880)
         );
  OAI222XL U1539 ( .A0(n911), .A1(n1460), .B0(n579), .B1(n1459), .C0(n912), 
        .C1(n1463), .Y(n879) );
  AOI222XL U1540 ( .A0(n883), .A1(n161), .B0(n160), .B1(n884), .C0(n126), .C1(
        n886), .Y(n882) );
  AO22X1 U1541 ( .A0(n552), .A1(n1529), .B0(sword[31]), .B1(n553), .Y(
        new_sword[31]) );
  OAI22XL U1542 ( .A0(sword[30]), .A1(n554), .B0(n555), .B1(n1527), .Y(n553)
         );
  OAI222XL U1543 ( .A0(n584), .A1(n1510), .B0(n1466), .B1(n1509), .C0(n585), 
        .C1(n1527), .Y(n552) );
  AOI222XL U1544 ( .A0(n556), .A1(n166), .B0(n165), .B1(n557), .C0(n136), .C1(
        n559), .Y(n555) );
  OA21XL U1545 ( .A0(n1157), .A1(n1158), .B0(n985), .Y(n1156) );
  OAI211X1 U1546 ( .A0(n1133), .A1(n32), .B0(n896), .C0(n1438), .Y(n1157) );
  OAI222XL U1547 ( .A0(n940), .A1(n1444), .B0(n992), .B1(n1428), .C0(sword[19]), .C1(n28), .Y(n1158) );
  OA21XL U1548 ( .A0(n836), .A1(n837), .B0(n689), .Y(n835) );
  OAI211X1 U1549 ( .A0(n812), .A1(n58), .B0(n569), .C0(n1489), .Y(n836) );
  OAI222XL U1550 ( .A0(n613), .A1(n1495), .B0(n696), .B1(n1479), .C0(sword[27]), .C1(n54), .Y(n837) );
  OA21XL U1551 ( .A0(n1070), .A1(n1071), .B0(n442), .Y(n1069) );
  OAI211X1 U1552 ( .A0(n666), .A1(n45), .B0(n353), .C0(n1513), .Y(n1070) );
  OAI222XL U1553 ( .A0(n397), .A1(n1519), .B0(n449), .B1(n182), .C0(sword[3]), 
        .C1(n11), .Y(n1071) );
  OA21XL U1554 ( .A0(n244), .A1(n245), .B0(n246), .Y(n243) );
  OAI211X1 U1555 ( .A0(n1548), .A1(n247), .B0(n204), .C0(n213), .Y(n245) );
  OAI222XL U1556 ( .A0(n144), .A1(sword[11]), .B0(n1545), .B1(n248), .C0(n194), 
        .C1(n249), .Y(n244) );
  OAI221XL U1557 ( .A0(n96), .A1(n18), .B0(n226), .B1(n148), .C0(n1266), .Y(
        n1264) );
  AOI2BB2X1 U1558 ( .B0(n1547), .B1(n289), .A0N(n146), .A1N(sword[10]), .Y(
        n1266) );
  NOR2X1 U1559 ( .A(sword[14]), .B(n97), .Y(n1274) );
  NOR2X1 U1560 ( .A(n1463), .B(sword[23]), .Y(n936) );
  NOR2X1 U1561 ( .A(n1541), .B(sword[7]), .Y(n393) );
  NOR2X1 U1562 ( .A(n1527), .B(sword[31]), .Y(n609) );
  NOR2X1 U1563 ( .A(sword[22]), .B(sword[23]), .Y(n1009) );
  NOR2X1 U1564 ( .A(sword[6]), .B(sword[7]), .Y(n466) );
  NOR2X1 U1565 ( .A(sword[30]), .B(sword[31]), .Y(n713) );
  NAND2X1 U1566 ( .A(sword[14]), .B(n97), .Y(n236) );
  BUFX2 U1567 ( .A(sword[15]), .Y(n97) );
  NAND2X1 U1568 ( .A(sword[23]), .B(sword[22]), .Y(n1122) );
  NAND2X1 U1569 ( .A(sword[31]), .B(sword[30]), .Y(n801) );
  NAND2X1 U1570 ( .A(sword[7]), .B(sword[6]), .Y(n655) );
  NAND2X1 U1571 ( .A(sword[23]), .B(n1463), .Y(n1120) );
  NAND2X1 U1572 ( .A(sword[31]), .B(n1527), .Y(n799) );
  NAND2X1 U1573 ( .A(sword[7]), .B(n1541), .Y(n653) );
  INVX1 U1574 ( .A(sword[23]), .Y(n1465) );
  INVX1 U1575 ( .A(sword[7]), .Y(n1543) );
  INVX1 U1576 ( .A(sword[31]), .Y(n1529) );
  INVX1 U1577 ( .A(sword[5]), .Y(n153) );
  INVX1 U1578 ( .A(sword[29]), .Y(n168) );
  INVX1 U1579 ( .A(sword[21]), .Y(n163) );
  INVX1 U1580 ( .A(sword[13]), .Y(n158) );
endmodule


module aes_decipher_block ( clk, reset_n, next, keylen, round, round_key, 
        block, new_block, ready );
  output [3:0] round;
  input [127:0] round_key;
  input [127:0] block;
  output [127:0] new_block;
  input clk, reset_n, next, keylen;
  output ready;
  wire   \dec_ctrl_reg[0] , n7, n8, n11, n13, n16, n20, n21, n22, n23, n24,
         n26, n27, n28, n29, n31, n32, n34, n35, n37, n38, n39, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n62, n63, n65, n67, n68, n69, n70, n71, n73, n76, n79, n80, n81,
         n83, n84, n86, n87, n89, n90, n92, n93, n94, n95, n98, n99, n100,
         n102, n103, n104, n105, n106, n109, n110, n112, n114, n117, n118,
         n119, n121, n122, n123, n124, n125, n126, n127, n129, n130, n132,
         n134, n136, n137, n138, n139, n140, n141, n142, n143, n145, n146,
         n148, n149, n150, n151, n152, n154, n157, n158, n159, n161, n163,
         n164, n167, n168, n169, n173, n175, n176, n177, n178, n179, n181,
         n182, n183, n184, n185, n186, n187, n188, n191, n193, n195, n196,
         n197, n198, n199, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1, n2, n3, n4, n5, n6, n9, n10, n12, n14,
         n15, n17, n18, n19, n25, n30, n33, n36, n40, n59, n60, n61, n64, n66,
         n72, n74, n75, n77, n78, n82, n85, n88, n91, n96, n97, n101, n107,
         n108, n111, n113, n115, n116, n120, n128, n131, n133, n135, n144,
         n147, n153, n155, n156, n160, n162, n165, n166, n170, n171, n172,
         n174, n180, n189, n190, n192, n194, n200, n239, n743, n1486, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710;
  wire   [31:0] tmp_sboxw;
  wire   [31:0] new_sboxw;
  wire   [1:0] sword_ctr_reg;

  aes_inv_sbox inv_sbox_inst ( .sword(tmp_sboxw), .new_sword(new_sboxw) );
  DFFSX1 ready_reg_reg ( .D(n1619), .CK(clk), .SN(n1652), .Q(ready) );
  DFFRX1 \block_w0_reg_reg[21]  ( .D(n1501), .CK(clk), .RN(n1647), .Q(
        new_block[117]), .QN(n169) );
  DFFRX1 \block_w0_reg_reg[29]  ( .D(n1493), .CK(clk), .RN(n1654), .Q(
        new_block[125]), .QN(n157) );
  DFFRX1 \block_w3_reg_reg[13]  ( .D(n1604), .CK(clk), .RN(n1643), .Q(
        new_block[13]), .QN(n39) );
  DFFRX1 \block_w3_reg_reg[5]  ( .D(n1612), .CK(clk), .RN(n1649), .Q(
        new_block[5]), .QN(n48) );
  DFFRX1 \block_w1_reg_reg[29]  ( .D(n1524), .CK(clk), .RN(n1648), .Q(
        new_block[93]), .QN(n112) );
  DFFRX1 \block_w1_reg_reg[21]  ( .D(n1532), .CK(clk), .RN(n1641), .Q(
        new_block[85]), .QN(n124) );
  DFFRX1 \block_w2_reg_reg[5]  ( .D(n1580), .CK(clk), .RN(n1647), .Q(
        new_block[37]), .QN(n100) );
  DFFRX1 \block_w2_reg_reg[29]  ( .D(n1556), .CK(clk), .RN(n1640), .Q(
        new_block[61]), .QN(n63) );
  DFFRX1 \block_w3_reg_reg[23]  ( .D(n1594), .CK(clk), .RN(n1647), .Q(
        new_block[23]), .QN(n26) );
  DFFRX1 \block_w3_reg_reg[22]  ( .D(n1595), .CK(clk), .RN(n1647), .Q(
        new_block[22]), .QN(n27) );
  DFFRX1 \block_w2_reg_reg[31]  ( .D(n1554), .CK(clk), .RN(n1648), .Q(
        new_block[63]), .QN(n58) );
  DFFRX1 \block_w0_reg_reg[15]  ( .D(n1507), .CK(clk), .RN(n1648), .Q(
        new_block[111]), .QN(n179) );
  DFFRX1 \block_w2_reg_reg[6]  ( .D(n1579), .CK(clk), .RN(n1649), .Q(
        new_block[38]), .QN(n99) );
  DFFRX1 \block_w3_reg_reg[14]  ( .D(n1603), .CK(clk), .RN(n1652), .Q(
        new_block[14]), .QN(n38) );
  DFFRX1 \block_w0_reg_reg[22]  ( .D(n1500), .CK(clk), .RN(n1651), .Q(
        new_block[118]), .QN(n168) );
  DFFRX1 \block_w2_reg_reg[14]  ( .D(n1571), .CK(clk), .RN(n1652), .Q(
        new_block[46]), .QN(n87) );
  DFFRX1 \block_w1_reg_reg[6]  ( .D(n1547), .CK(clk), .RN(n1653), .Q(
        new_block[70]), .QN(n143) );
  DFFRX1 \block_w0_reg_reg[13]  ( .D(n1509), .CK(clk), .RN(n1651), .Q(
        new_block[109]), .QN(n182) );
  DFFRX1 \block_w1_reg_reg[7]  ( .D(n1546), .CK(clk), .RN(n1650), .Q(
        new_block[71]), .QN(n142) );
  DFFRX1 \block_w0_reg_reg[7]  ( .D(n1515), .CK(clk), .RN(n1650), .Q(
        new_block[103]), .QN(n188) );
  DFFRX1 \block_w1_reg_reg[30]  ( .D(n1523), .CK(clk), .RN(n1641), .Q(
        new_block[94]), .QN(n110) );
  DFFRX1 \block_w3_reg_reg[7]  ( .D(n1610), .CK(clk), .RN(n1640), .Q(
        new_block[7]), .QN(n46) );
  DFFRX1 \block_w0_reg_reg[30]  ( .D(n1492), .CK(clk), .RN(n1652), .Q(
        new_block[126]), .QN(n154) );
  DFFRX1 \block_w0_reg_reg[31]  ( .D(n1491), .CK(clk), .RN(n1651), .Q(
        new_block[127]), .QN(n152) );
  DFFRX1 \block_w3_reg_reg[21]  ( .D(n1596), .CK(clk), .RN(n1646), .Q(
        new_block[21]), .QN(n28) );
  DFFRX1 \block_w3_reg_reg[6]  ( .D(n1611), .CK(clk), .RN(n1651), .Q(
        new_block[6]), .QN(n47) );
  DFFRX1 \block_w0_reg_reg[14]  ( .D(n1508), .CK(clk), .RN(n1654), .Q(
        new_block[110]), .QN(n181) );
  DFFRX1 \block_w0_reg_reg[5]  ( .D(n1517), .CK(clk), .RN(n1641), .Q(
        new_block[101]), .QN(n193) );
  DFFRX1 \block_w0_reg_reg[6]  ( .D(n1516), .CK(clk), .RN(n1640), .Q(
        new_block[102]), .QN(n191) );
  DFFRX1 \block_w0_reg_reg[23]  ( .D(n1499), .CK(clk), .RN(n1641), .Q(
        new_block[119]), .QN(n167) );
  DFFRX1 \block_w3_reg_reg[29]  ( .D(n1588), .CK(clk), .RN(n1643), .Q(
        new_block[29]), .QN(n16) );
  DFFRX1 \block_w3_reg_reg[30]  ( .D(n1587), .CK(clk), .RN(n1644), .Q(
        new_block[30]), .QN(n13) );
  DFFRX1 \block_w3_reg_reg[31]  ( .D(n1586), .CK(clk), .RN(n1645), .Q(
        new_block[31]), .QN(n11) );
  DFFRX1 \block_w3_reg_reg[15]  ( .D(n1602), .CK(clk), .RN(n1649), .Q(
        new_block[15]), .QN(n37) );
  DFFRX1 \block_w1_reg_reg[22]  ( .D(n1531), .CK(clk), .RN(n1650), .Q(
        new_block[86]), .QN(n123) );
  DFFRX1 \block_w1_reg_reg[31]  ( .D(n1522), .CK(clk), .RN(n1650), .Q(
        new_block[95]), .QN(n109) );
  DFFRX1 \block_w1_reg_reg[23]  ( .D(n1530), .CK(clk), .RN(n1650), .Q(
        new_block[87]), .QN(n122) );
  DFFRX1 \block_w2_reg_reg[30]  ( .D(n1555), .CK(clk), .RN(n1654), .Q(
        new_block[62]), .QN(n62) );
  DFFRX1 \block_w2_reg_reg[23]  ( .D(n1562), .CK(clk), .RN(n1650), .Q(
        new_block[55]), .QN(n71) );
  DFFRX1 \block_w1_reg_reg[13]  ( .D(n1540), .CK(clk), .RN(n1644), .Q(
        new_block[77]), .QN(n136) );
  DFFRX1 \block_w1_reg_reg[5]  ( .D(n1548), .CK(clk), .RN(n1644), .Q(
        new_block[69]), .QN(n145) );
  DFFRX1 \block_w1_reg_reg[14]  ( .D(n1539), .CK(clk), .RN(n1645), .Q(
        new_block[78]), .QN(n134) );
  DFFRX1 \block_w1_reg_reg[15]  ( .D(n1538), .CK(clk), .RN(n1652), .Q(
        new_block[79]), .QN(n132) );
  DFFRX1 \block_w2_reg_reg[13]  ( .D(n1572), .CK(clk), .RN(n1647), .Q(
        new_block[45]), .QN(n89) );
  DFFRX1 \block_w2_reg_reg[7]  ( .D(n1578), .CK(clk), .RN(n1652), .Q(
        new_block[39]), .QN(n98) );
  DFFRX1 \block_w2_reg_reg[22]  ( .D(n1563), .CK(clk), .RN(n1651), .Q(
        new_block[54]), .QN(n73) );
  DFFRX1 \block_w2_reg_reg[15]  ( .D(n1570), .CK(clk), .RN(n1640), .Q(
        new_block[47]), .QN(n86) );
  DFFRX1 \block_w2_reg_reg[21]  ( .D(n1564), .CK(clk), .RN(n1651), .Q(
        new_block[53]), .QN(n76) );
  DFFRX1 \block_w0_reg_reg[0]  ( .D(n1618), .CK(clk), .RN(n1642), .Q(
        new_block[96]), .QN(n199) );
  DFFRX1 \block_w0_reg_reg[2]  ( .D(n1520), .CK(clk), .RN(n1646), .Q(
        new_block[98]), .QN(n197) );
  DFFRX1 \block_w0_reg_reg[17]  ( .D(n1505), .CK(clk), .RN(n1647), .Q(
        new_block[113]), .QN(n177) );
  DFFRX1 \block_w0_reg_reg[18]  ( .D(n1504), .CK(clk), .RN(n1648), .Q(
        new_block[114]), .QN(n176) );
  DFFRX1 \block_w0_reg_reg[16]  ( .D(n1506), .CK(clk), .RN(n1649), .Q(
        new_block[112]), .QN(n178) );
  DFFRX1 \block_w0_reg_reg[24]  ( .D(n1498), .CK(clk), .RN(n1649), .Q(
        new_block[120]), .QN(n164) );
  DFFRX1 \block_w0_reg_reg[3]  ( .D(n1519), .CK(clk), .RN(n1649), .Q(
        new_block[99]), .QN(n196) );
  DFFRX1 \block_w0_reg_reg[11]  ( .D(n1511), .CK(clk), .RN(n1654), .Q(
        new_block[107]), .QN(n184) );
  DFFRX1 \block_w0_reg_reg[9]  ( .D(n1513), .CK(clk), .RN(n1653), .Q(
        new_block[105]), .QN(n186) );
  DFFRX1 \block_w0_reg_reg[12]  ( .D(n1510), .CK(clk), .RN(n1641), .Q(
        new_block[108]), .QN(n183) );
  DFFRX1 \block_w0_reg_reg[8]  ( .D(n1514), .CK(clk), .RN(n1653), .Q(
        new_block[104]), .QN(n187) );
  DFFRX1 \block_w3_reg_reg[1]  ( .D(n1616), .CK(clk), .RN(n1642), .Q(
        new_block[1]), .QN(n52) );
  DFFRX1 \block_w3_reg_reg[26]  ( .D(n1591), .CK(clk), .RN(n1643), .Q(
        new_block[26]), .QN(n22) );
  DFFRX1 \block_w3_reg_reg[27]  ( .D(n1590), .CK(clk), .RN(n1643), .Q(
        new_block[27]), .QN(n21) );
  DFFRX1 \block_w3_reg_reg[19]  ( .D(n1598), .CK(clk), .RN(n1644), .Q(
        new_block[19]), .QN(n31) );
  DFFRX1 \block_w3_reg_reg[11]  ( .D(n1606), .CK(clk), .RN(n1644), .Q(
        new_block[11]), .QN(n42) );
  DFFRX1 \block_w3_reg_reg[18]  ( .D(n1599), .CK(clk), .RN(n1645), .Q(
        new_block[18]), .QN(n32) );
  DFFRX1 \block_w3_reg_reg[24]  ( .D(n1593), .CK(clk), .RN(n1646), .Q(
        new_block[24]), .QN(n24) );
  DFFRX1 \block_w3_reg_reg[16]  ( .D(n1601), .CK(clk), .RN(n1646), .Q(
        new_block[16]), .QN(n35) );
  DFFRX1 \block_w3_reg_reg[4]  ( .D(n1613), .CK(clk), .RN(n1646), .Q(
        new_block[4]), .QN(n49) );
  DFFRX1 \block_w3_reg_reg[8]  ( .D(n1609), .CK(clk), .RN(n1647), .Q(
        new_block[8]), .QN(n45) );
  DFFRX1 \block_w3_reg_reg[2]  ( .D(n1615), .CK(clk), .RN(n1648), .Q(
        new_block[2]), .QN(n51) );
  DFFRX1 \block_w1_reg_reg[9]  ( .D(n1544), .CK(clk), .RN(n1643), .Q(
        new_block[73]), .QN(n140) );
  DFFRX1 \block_w1_reg_reg[10]  ( .D(n1543), .CK(clk), .RN(n1644), .Q(
        new_block[74]), .QN(n139) );
  DFFRX1 \block_w1_reg_reg[11]  ( .D(n1542), .CK(clk), .RN(n1645), .Q(
        new_block[75]), .QN(n138) );
  DFFRX1 \block_w1_reg_reg[8]  ( .D(n1545), .CK(clk), .RN(n1646), .Q(
        new_block[72]), .QN(n141) );
  DFFRX1 \block_w1_reg_reg[26]  ( .D(n1527), .CK(clk), .RN(n1646), .Q(
        new_block[90]), .QN(n118) );
  DFFRX1 \block_w1_reg_reg[28]  ( .D(n1525), .CK(clk), .RN(n1654), .Q(
        new_block[92]), .QN(n114) );
  DFFRX1 \block_w1_reg_reg[18]  ( .D(n1535), .CK(clk), .RN(n1650), .Q(
        new_block[82]), .QN(n127) );
  DFFRX1 \block_w1_reg_reg[27]  ( .D(n1526), .CK(clk), .RN(n1650), .Q(
        new_block[91]), .QN(n117) );
  DFFRX1 \block_w1_reg_reg[20]  ( .D(n1533), .CK(clk), .RN(n1654), .Q(
        new_block[84]), .QN(n125) );
  DFFRX1 \block_w1_reg_reg[16]  ( .D(n1537), .CK(clk), .RN(n1652), .Q(
        new_block[80]), .QN(n130) );
  DFFRX1 \block_w1_reg_reg[25]  ( .D(n1528), .CK(clk), .RN(n1641), .Q(
        new_block[89]), .QN(n119) );
  DFFRX1 \block_w2_reg_reg[3]  ( .D(n1582), .CK(clk), .RN(n1643), .Q(
        new_block[35]), .QN(n103) );
  DFFRX1 \block_w2_reg_reg[18]  ( .D(n1567), .CK(clk), .RN(n1645), .Q(
        new_block[50]), .QN(n81) );
  DFFRX1 \block_w2_reg_reg[0]  ( .D(n1585), .CK(clk), .RN(n1646), .Q(
        new_block[32]), .QN(n106) );
  DFFRX1 \block_w2_reg_reg[2]  ( .D(n1583), .CK(clk), .RN(n1646), .Q(
        new_block[34]), .QN(n104) );
  DFFRX1 \block_w2_reg_reg[25]  ( .D(n1560), .CK(clk), .RN(n1648), .Q(
        new_block[57]), .QN(n69) );
  DFFRX1 \block_w2_reg_reg[28]  ( .D(n1557), .CK(clk), .RN(n1648), .Q(
        new_block[60]), .QN(n65) );
  DFFRX1 \block_w2_reg_reg[19]  ( .D(n1566), .CK(clk), .RN(n1649), .Q(
        new_block[51]), .QN(n80) );
  DFFRX1 \block_w2_reg_reg[8]  ( .D(n1577), .CK(clk), .RN(n1652), .Q(
        new_block[40]), .QN(n95) );
  DFFRX1 \block_w2_reg_reg[24]  ( .D(n1561), .CK(clk), .RN(n1651), .Q(
        new_block[56]), .QN(n70) );
  DFFRX1 \block_w0_reg_reg[27]  ( .D(n1495), .CK(clk), .RN(n1654), .Q(
        new_block[123]), .QN(n159) );
  DFFRX1 \block_w0_reg_reg[10]  ( .D(n1512), .CK(clk), .RN(n1651), .Q(
        new_block[106]), .QN(n185) );
  DFFRX1 \block_w0_reg_reg[28]  ( .D(n1494), .CK(clk), .RN(n1641), .Q(
        new_block[124]), .QN(n158) );
  DFFRX1 \block_w0_reg_reg[1]  ( .D(n1521), .CK(clk), .RN(n1640), .Q(
        new_block[97]), .QN(n198) );
  DFFRX1 \block_w0_reg_reg[26]  ( .D(n1496), .CK(clk), .RN(n1641), .Q(
        new_block[122]), .QN(n161) );
  DFFRX1 \block_w3_reg_reg[25]  ( .D(n1592), .CK(clk), .RN(n1643), .Q(
        new_block[25]), .QN(n23) );
  DFFRX1 \block_w3_reg_reg[10]  ( .D(n1607), .CK(clk), .RN(n1643), .Q(
        new_block[10]), .QN(n43) );
  DFFRX1 \block_w3_reg_reg[9]  ( .D(n1608), .CK(clk), .RN(n1644), .Q(
        new_block[9]), .QN(n44) );
  DFFRX1 \block_w3_reg_reg[3]  ( .D(n1614), .CK(clk), .RN(n1645), .Q(
        new_block[3]), .QN(n50) );
  DFFRX1 \block_w3_reg_reg[20]  ( .D(n1597), .CK(clk), .RN(n1645), .Q(
        new_block[20]), .QN(n29) );
  DFFRX1 \block_w3_reg_reg[0]  ( .D(n1617), .CK(clk), .RN(n1640), .Q(
        new_block[0]), .QN(n53) );
  DFFRX1 \block_w0_reg_reg[19]  ( .D(n1503), .CK(clk), .RN(n1645), .Q(
        new_block[115]), .QN(n175) );
  DFFRX1 \block_w0_reg_reg[25]  ( .D(n1497), .CK(clk), .RN(n1647), .Q(
        new_block[121]), .QN(n163) );
  DFFRX1 \block_w0_reg_reg[20]  ( .D(n1502), .CK(clk), .RN(n1648), .Q(
        new_block[116]), .QN(n173) );
  DFFRX1 \block_w0_reg_reg[4]  ( .D(n1518), .CK(clk), .RN(n1650), .Q(
        new_block[100]), .QN(n195) );
  DFFRX1 \block_w3_reg_reg[28]  ( .D(n1589), .CK(clk), .RN(n1643), .Q(
        new_block[28]), .QN(n20) );
  DFFRX1 \block_w3_reg_reg[17]  ( .D(n1600), .CK(clk), .RN(n1644), .Q(
        new_block[17]), .QN(n34) );
  DFFRX1 \block_w3_reg_reg[12]  ( .D(n1605), .CK(clk), .RN(n1645), .Q(
        new_block[12]), .QN(n41) );
  DFFRX1 \block_w1_reg_reg[12]  ( .D(n1541), .CK(clk), .RN(n1643), .Q(
        new_block[76]), .QN(n137) );
  DFFRX1 \block_w1_reg_reg[0]  ( .D(n1553), .CK(clk), .RN(n1647), .Q(
        new_block[64]), .QN(n151) );
  DFFRX1 \block_w1_reg_reg[2]  ( .D(n1551), .CK(clk), .RN(n1648), .Q(
        new_block[66]), .QN(n149) );
  DFFRX1 \block_w1_reg_reg[4]  ( .D(n1549), .CK(clk), .RN(n1649), .Q(
        new_block[68]), .QN(n146) );
  DFFRX1 \block_w1_reg_reg[19]  ( .D(n1534), .CK(clk), .RN(n1649), .Q(
        new_block[83]), .QN(n126) );
  DFFRX1 \block_w1_reg_reg[1]  ( .D(n1552), .CK(clk), .RN(n1654), .Q(
        new_block[65]), .QN(n150) );
  DFFRX1 \block_w2_reg_reg[1]  ( .D(n1584), .CK(clk), .RN(n1644), .Q(
        new_block[33]), .QN(n105) );
  DFFRX1 \block_w2_reg_reg[16]  ( .D(n1569), .CK(clk), .RN(n1645), .Q(
        new_block[48]), .QN(n84) );
  DFFRX1 \block_w2_reg_reg[26]  ( .D(n1559), .CK(clk), .RN(n1646), .Q(
        new_block[58]), .QN(n68) );
  DFFRX1 \block_w2_reg_reg[10]  ( .D(n1575), .CK(clk), .RN(n1648), .Q(
        new_block[42]), .QN(n93) );
  DFFRX1 \block_w2_reg_reg[27]  ( .D(n1558), .CK(clk), .RN(n1649), .Q(
        new_block[59]), .QN(n67) );
  DFFRX1 \block_w2_reg_reg[12]  ( .D(n1573), .CK(clk), .RN(n1653), .Q(
        new_block[44]), .QN(n90) );
  DFFRX1 \block_w2_reg_reg[9]  ( .D(n1576), .CK(clk), .RN(n1641), .Q(
        new_block[41]), .QN(n94) );
  DFFRX1 \block_w1_reg_reg[3]  ( .D(n1550), .CK(clk), .RN(n1653), .Q(
        new_block[67]), .QN(n148) );
  DFFRX1 \block_w1_reg_reg[24]  ( .D(n1529), .CK(clk), .RN(n1653), .Q(
        new_block[88]), .QN(n121) );
  DFFRX1 \block_w1_reg_reg[17]  ( .D(n1536), .CK(clk), .RN(n1640), .Q(
        new_block[81]), .QN(n129) );
  DFFRX1 \block_w2_reg_reg[4]  ( .D(n1581), .CK(clk), .RN(n1644), .Q(
        new_block[36]), .QN(n102) );
  DFFRX1 \block_w2_reg_reg[11]  ( .D(n1574), .CK(clk), .RN(n1647), .Q(
        new_block[43]), .QN(n92) );
  DFFRX1 \block_w2_reg_reg[17]  ( .D(n1568), .CK(clk), .RN(n1653), .Q(
        new_block[49]), .QN(n83) );
  DFFRX1 \block_w2_reg_reg[20]  ( .D(n1565), .CK(clk), .RN(n1650), .Q(
        new_block[52]), .QN(n79) );
  DFFRX1 \sword_ctr_reg_reg[1]  ( .D(n1626), .CK(clk), .RN(n1642), .Q(
        sword_ctr_reg[1]), .QN(n56) );
  DFFRX1 \sword_ctr_reg_reg[0]  ( .D(n1627), .CK(clk), .RN(n1642), .Q(
        sword_ctr_reg[0]), .QN(n57) );
  DFFRX1 \round_ctr_reg_reg[1]  ( .D(n1622), .CK(clk), .RN(n1642), .Q(round[1]), .QN(n54) );
  DFFRX1 \round_ctr_reg_reg[0]  ( .D(n1623), .CK(clk), .RN(n1642), .Q(round[0]), .QN(n55) );
  DFFRX1 \round_ctr_reg_reg[3]  ( .D(n1620), .CK(clk), .RN(n1642), .Q(round[3]) );
  DFFRX1 \round_ctr_reg_reg[2]  ( .D(n1621), .CK(clk), .RN(n1642), .Q(round[2]) );
  DFFRX1 \dec_ctrl_reg_reg[0]  ( .D(n1624), .CK(clk), .RN(n1642), .Q(
        \dec_ctrl_reg[0] ), .QN(n8) );
  DFFRX1 \dec_ctrl_reg_reg[1]  ( .D(n1625), .CK(clk), .RN(n1642), .Q(n1), .QN(
        n7) );
  OAI221XL U3 ( .A0(n1637), .A1(n41), .B0(n1634), .B1(n183), .C0(n233), .Y(
        tmp_sboxw[12]) );
  OAI221XL U4 ( .A0(n1637), .A1(n42), .B0(n1634), .B1(n184), .C0(n234), .Y(
        tmp_sboxw[11]) );
  OAI221XL U5 ( .A0(n1638), .A1(n50), .B0(n1636), .B1(n196), .C0(n211), .Y(
        tmp_sboxw[3]) );
  OAI221XL U6 ( .A0(n1638), .A1(n49), .B0(n1636), .B1(n195), .C0(n210), .Y(
        tmp_sboxw[4]) );
  OAI221XL U7 ( .A0(n1638), .A1(n21), .B0(n1636), .B1(n159), .C0(n217), .Y(
        tmp_sboxw[27]) );
  OAI221XL U8 ( .A0(n1638), .A1(n20), .B0(n1636), .B1(n158), .C0(n216), .Y(
        tmp_sboxw[28]) );
  OAI221XL U9 ( .A0(n1639), .A1(n31), .B0(n1635), .B1(n175), .C0(n226), .Y(
        tmp_sboxw[19]) );
  OAI221XL U10 ( .A0(n1639), .A1(n29), .B0(n1635), .B1(n173), .C0(n224), .Y(
        tmp_sboxw[20]) );
  OAI221XL U11 ( .A0(n1637), .A1(n38), .B0(n1634), .B1(n181), .C0(n231), .Y(
        tmp_sboxw[14]) );
  NAND2X1 U12 ( .A(n861), .B(n1634), .Y(n2) );
  NAND2X1 U13 ( .A(n1474), .B(n1704), .Y(n238) );
  NOR2X1 U14 ( .A(n1475), .B(n1474), .Y(n244) );
  XOR2X1 U15 ( .A(new_block[7]), .B(round_key[7]), .Y(n777) );
  XOR2X1 U16 ( .A(new_block[23]), .B(round_key[23]), .Y(n710) );
  XOR2X1 U17 ( .A(new_block[71]), .B(round_key[71]), .Y(n567) );
  XOR2X1 U18 ( .A(new_block[63]), .B(round_key[63]), .Y(n859) );
  OAI221XL U19 ( .A0(n1639), .A1(n44), .B0(n202), .B1(n186), .C0(n203), .Y(
        tmp_sboxw[9]) );
  OAI221XL U20 ( .A0(n1639), .A1(n45), .B0(n202), .B1(n187), .C0(n206), .Y(
        tmp_sboxw[8]) );
  OAI221XL U21 ( .A0(n1639), .A1(n23), .B0(n1635), .B1(n163), .C0(n219), .Y(
        tmp_sboxw[25]) );
  OAI221XL U22 ( .A0(n1639), .A1(n24), .B0(n1635), .B1(n164), .C0(n220), .Y(
        tmp_sboxw[24]) );
  OAI221XL U23 ( .A0(n1639), .A1(n52), .B0(n1635), .B1(n198), .C0(n225), .Y(
        tmp_sboxw[1]) );
  XOR2X1 U24 ( .A(n86), .B(round_key[47]), .Y(n1236) );
  XOR2X1 U25 ( .A(n132), .B(round_key[79]), .Y(n1358) );
  NOR2X1 U26 ( .A(n7), .B(\dec_ctrl_reg[0] ), .Y(n1489) );
  OAI221XL U27 ( .A0(n1637), .A1(n35), .B0(n1634), .B1(n178), .C0(n229), .Y(
        tmp_sboxw[16]) );
  OAI221XL U28 ( .A0(n1637), .A1(n53), .B0(n1634), .B1(n199), .C0(n236), .Y(
        tmp_sboxw[0]) );
  OAI221XL U29 ( .A0(n1637), .A1(n34), .B0(n1634), .B1(n177), .C0(n228), .Y(
        tmp_sboxw[17]) );
  XOR2X1 U30 ( .A(new_block[126]), .B(round_key[126]), .Y(n251) );
  XNOR2X1 U31 ( .A(n47), .B(round_key[6]), .Y(n338) );
  XNOR2X1 U32 ( .A(n62), .B(round_key[62]), .Y(n417) );
  XOR2X1 U33 ( .A(new_block[118]), .B(round_key[118]), .Y(n333) );
  XOR2X1 U34 ( .A(new_block[46]), .B(round_key[46]), .Y(n879) );
  XOR2X1 U35 ( .A(new_block[22]), .B(round_key[22]), .Y(n1088) );
  XOR2X1 U36 ( .A(new_block[111]), .B(round_key[111]), .Y(n404) );
  XOR2X1 U37 ( .A(new_block[38]), .B(round_key[38]), .Y(n785) );
  XOR2X1 U38 ( .A(new_block[14]), .B(round_key[14]), .Y(n712) );
  XOR2X1 U39 ( .A(new_block[103]), .B(round_key[103]), .Y(n484) );
  XOR2X1 U40 ( .A(new_block[94]), .B(round_key[94]), .Y(n569) );
  XOR2X1 U41 ( .A(new_block[127]), .B(round_key[127]), .Y(n243) );
  XOR2X1 U42 ( .A(n181), .B(round_key[110]), .Y(n641) );
  XOR2X1 U43 ( .A(n134), .B(round_key[78]), .Y(n577) );
  XOR2X1 U44 ( .A(n13), .B(round_key[30]), .Y(n720) );
  XOR2X1 U45 ( .A(n76), .B(round_key[53]), .Y(n877) );
  XOR2X1 U46 ( .A(n83), .B(round_key[49]), .Y(n927) );
  OAI221XL U47 ( .A0(n1637), .A1(n37), .B0(n1634), .B1(n179), .C0(n230), .Y(
        tmp_sboxw[15]) );
  BUFX2 U48 ( .A(n1653), .Y(n1650) );
  BUFX2 U49 ( .A(n1651), .Y(n1649) );
  BUFX2 U50 ( .A(n1651), .Y(n1648) );
  BUFX2 U51 ( .A(n1652), .Y(n1647) );
  BUFX2 U52 ( .A(n1652), .Y(n1646) );
  BUFX2 U53 ( .A(n1653), .Y(n1645) );
  BUFX2 U54 ( .A(n1653), .Y(n1644) );
  BUFX2 U55 ( .A(n1654), .Y(n1643) );
  BUFX2 U56 ( .A(n1654), .Y(n1642) );
  BUFX2 U57 ( .A(n1640), .Y(n1651) );
  BUFX2 U58 ( .A(n1640), .Y(n1652) );
  BUFX2 U59 ( .A(n1640), .Y(n1653) );
  BUFX2 U60 ( .A(reset_n), .Y(n1640) );
  BUFX2 U61 ( .A(n1641), .Y(n1654) );
  BUFX2 U62 ( .A(reset_n), .Y(n1641) );
  BUFX2 U63 ( .A(n559), .Y(n40) );
  BUFX2 U64 ( .A(n864), .Y(n18) );
  BUFX2 U65 ( .A(n1150), .Y(n9) );
  BUFX2 U66 ( .A(n165), .Y(n160) );
  BUFX2 U67 ( .A(n241), .Y(n156) );
  BUFX2 U68 ( .A(n241), .Y(n155) );
  BUFX2 U69 ( .A(n241), .Y(n153) );
  BUFX2 U70 ( .A(n561), .Y(n30) );
  BUFX2 U71 ( .A(n561), .Y(n33) );
  BUFX2 U72 ( .A(n866), .Y(n17) );
  BUFX2 U73 ( .A(n866), .Y(n15) );
  BUFX2 U74 ( .A(n866), .Y(n14) );
  BUFX2 U75 ( .A(n1152), .Y(n5) );
  BUFX2 U76 ( .A(n1152), .Y(n6) );
  BUFX2 U77 ( .A(n1152), .Y(n4) );
  BUFX2 U78 ( .A(n561), .Y(n36) );
  BUFX2 U79 ( .A(n559), .Y(n60) );
  BUFX2 U80 ( .A(n864), .Y(n25) );
  BUFX2 U81 ( .A(n864), .Y(n19) );
  BUFX2 U82 ( .A(n1150), .Y(n10) );
  BUFX2 U83 ( .A(n559), .Y(n59) );
  BUFX2 U84 ( .A(n1150), .Y(n12) );
  BUFX2 U85 ( .A(n144), .Y(n115) );
  BUFX2 U86 ( .A(n133), .Y(n111) );
  BUFX2 U87 ( .A(n131), .Y(n120) );
  BUFX2 U88 ( .A(n144), .Y(n113) );
  BUFX2 U89 ( .A(n133), .Y(n116) );
  BUFX2 U90 ( .A(n131), .Y(n128) );
  BUFX2 U91 ( .A(n239), .Y(n172) );
  BUFX2 U92 ( .A(n200), .Y(n180) );
  BUFX2 U93 ( .A(n194), .Y(n190) );
  BUFX2 U94 ( .A(n200), .Y(n174) );
  BUFX2 U95 ( .A(n743), .Y(n166) );
  BUFX2 U96 ( .A(n194), .Y(n189) );
  BUFX2 U97 ( .A(n239), .Y(n171) );
  BUFX2 U98 ( .A(n743), .Y(n170) );
  BUFX2 U99 ( .A(n165), .Y(n162) );
  BUFX2 U100 ( .A(n200), .Y(n192) );
  XNOR2X1 U101 ( .A(n958), .B(n1323), .Y(n499) );
  XNOR2X1 U102 ( .A(n887), .B(n1245), .Y(n419) );
  XNOR2X1 U103 ( .A(n1096), .B(n1165), .Y(n339) );
  XOR2X1 U104 ( .A(n1026), .B(n1399), .Y(n259) );
  XOR2X1 U105 ( .A(n965), .B(n966), .Y(n516) );
  XOR2X1 U106 ( .A(n957), .B(n1323), .Y(n583) );
  XOR2X1 U107 ( .A(n886), .B(n1245), .Y(n800) );
  XOR2X1 U108 ( .A(n1025), .B(n1399), .Y(n656) );
  XOR2X1 U109 ( .A(n1095), .B(n1165), .Y(n726) );
  XNOR2X1 U110 ( .A(n817), .B(n818), .Y(n816) );
  XNOR2X1 U111 ( .A(n601), .B(n602), .Y(n600) );
  XOR2X1 U112 ( .A(n308), .B(n309), .Y(n307) );
  XOR2X1 U113 ( .A(n692), .B(n309), .Y(n1454) );
  XOR2X1 U114 ( .A(n388), .B(n1135), .Y(n1134) );
  XOR2X1 U115 ( .A(n762), .B(n1135), .Y(n1219) );
  XOR2X1 U116 ( .A(n976), .B(n602), .Y(n975) );
  XOR2X1 U117 ( .A(n529), .B(n527), .Y(n976) );
  XOR2X1 U118 ( .A(n904), .B(n818), .Y(n903) );
  XOR2X1 U119 ( .A(n448), .B(n446), .Y(n904) );
  INVX1 U120 ( .A(n831), .Y(n1673) );
  INVX1 U121 ( .A(n1129), .Y(n1687) );
  NOR3BXL U122 ( .AN(n238), .B(n244), .C(n108), .Y(n861) );
  NAND2X1 U123 ( .A(n861), .B(n1630), .Y(n864) );
  NAND2X1 U124 ( .A(n861), .B(n1631), .Y(n559) );
  NAND2X1 U125 ( .A(n861), .B(n1637), .Y(n1150) );
  AND2X2 U126 ( .A(n860), .B(n18), .Y(n866) );
  AND2X2 U127 ( .A(n860), .B(n40), .Y(n561) );
  AND2X2 U128 ( .A(n860), .B(n9), .Y(n1152) );
  AND2X2 U129 ( .A(n860), .B(n160), .Y(n241) );
  BUFX2 U130 ( .A(n2), .Y(n165) );
  BUFX2 U131 ( .A(n238), .Y(n1486) );
  BUFX2 U132 ( .A(n238), .Y(n200) );
  BUFX2 U133 ( .A(n238), .Y(n194) );
  BUFX2 U134 ( .A(n238), .Y(n239) );
  BUFX2 U135 ( .A(n238), .Y(n743) );
  BUFX2 U136 ( .A(n101), .Y(n135) );
  BUFX2 U137 ( .A(n135), .Y(n144) );
  BUFX2 U138 ( .A(n101), .Y(n133) );
  BUFX2 U139 ( .A(n101), .Y(n131) );
  BUFX2 U140 ( .A(n91), .Y(n72) );
  BUFX2 U141 ( .A(n88), .Y(n75) );
  BUFX2 U142 ( .A(n85), .Y(n78) );
  BUFX2 U143 ( .A(n88), .Y(n74) );
  BUFX2 U144 ( .A(n96), .Y(n61) );
  BUFX2 U145 ( .A(n85), .Y(n77) );
  BUFX2 U146 ( .A(n91), .Y(n66) );
  BUFX2 U147 ( .A(n96), .Y(n64) );
  BUFX2 U148 ( .A(n96), .Y(n82) );
  NOR2X1 U149 ( .A(n1704), .B(n1474), .Y(n860) );
  BUFX2 U150 ( .A(n204), .Y(n1631) );
  BUFX2 U151 ( .A(n204), .Y(n1632) );
  BUFX2 U152 ( .A(n204), .Y(n1633) );
  BUFX2 U153 ( .A(n205), .Y(n1628) );
  BUFX2 U154 ( .A(n205), .Y(n1629) );
  BUFX2 U155 ( .A(n201), .Y(n1637) );
  BUFX2 U156 ( .A(n201), .Y(n1638) );
  BUFX2 U157 ( .A(n205), .Y(n1630) );
  BUFX2 U158 ( .A(n201), .Y(n1639) );
  XNOR2X1 U159 ( .A(n1212), .B(n1136), .Y(n1129) );
  XOR2X1 U160 ( .A(n1447), .B(n1063), .Y(n692) );
  XOR2X1 U161 ( .A(n923), .B(n924), .Y(n468) );
  XOR2X1 U162 ( .A(n1365), .B(n997), .Y(n623) );
  XOR2X1 U163 ( .A(n1435), .B(n1422), .Y(n289) );
  XOR2X1 U164 ( .A(n1438), .B(n1439), .Y(n1435) );
  XNOR2X1 U165 ( .A(n1064), .B(n694), .Y(n1438) );
  XOR2X1 U166 ( .A(n1693), .B(n311), .Y(n1439) );
  XOR2X1 U167 ( .A(n1196), .B(n1184), .Y(n368) );
  XOR2X1 U168 ( .A(n1198), .B(n1199), .Y(n1196) );
  XNOR2X1 U169 ( .A(n393), .B(n764), .Y(n1198) );
  XOR2X1 U170 ( .A(n1200), .B(n390), .Y(n1199) );
  XOR2X1 U171 ( .A(n1276), .B(n1264), .Y(n448) );
  XOR2X1 U172 ( .A(n1279), .B(n1280), .Y(n1276) );
  XOR2X1 U173 ( .A(n1684), .B(n472), .Y(n1279) );
  XOR2X1 U174 ( .A(n844), .B(n926), .Y(n1280) );
  XOR2X1 U175 ( .A(n1365), .B(n996), .Y(n541) );
  XNOR2X1 U176 ( .A(n683), .B(n1440), .Y(n309) );
  XOR2X1 U177 ( .A(n955), .B(n956), .Y(n506) );
  XOR2X1 U178 ( .A(n957), .B(n958), .Y(n955) );
  XOR2X1 U179 ( .A(n1093), .B(n1094), .Y(n347) );
  XOR2X1 U180 ( .A(n1095), .B(n1096), .Y(n1093) );
  XOR2X1 U181 ( .A(n1656), .B(n249), .Y(n1072) );
  XOR2X1 U182 ( .A(n1690), .B(n328), .Y(n1144) );
  XNOR2X1 U183 ( .A(n624), .B(n557), .Y(n540) );
  XOR2X1 U184 ( .A(n1023), .B(n1024), .Y(n267) );
  XOR2X1 U185 ( .A(n1025), .B(n1026), .Y(n1023) );
  XOR2X1 U186 ( .A(n1677), .B(n409), .Y(n855) );
  XOR2X1 U187 ( .A(n1669), .B(n489), .Y(n1385) );
  XOR2X1 U188 ( .A(n390), .B(n764), .Y(n382) );
  XOR2X1 U189 ( .A(n472), .B(n844), .Y(n460) );
  XOR2X1 U190 ( .A(n469), .B(n926), .Y(n830) );
  XNOR2X1 U191 ( .A(n1188), .B(n1187), .Y(n745) );
  XOR2X1 U192 ( .A(n1037), .B(n318), .Y(n649) );
  XOR2X1 U193 ( .A(n898), .B(n480), .Y(n792) );
  XNOR2X1 U194 ( .A(n1330), .B(n1320), .Y(n966) );
  XNOR2X1 U195 ( .A(n977), .B(n532), .Y(n1330) );
  XNOR2X1 U196 ( .A(n1046), .B(n1047), .Y(n287) );
  XOR2X1 U197 ( .A(n1037), .B(n667), .Y(n643) );
  XOR2X1 U198 ( .A(n898), .B(n811), .Y(n870) );
  XOR2X1 U199 ( .A(n1107), .B(n737), .Y(n1079) );
  XOR2X1 U200 ( .A(n969), .B(n593), .Y(n942) );
  XNOR2X1 U201 ( .A(n1344), .B(n1343), .Y(n601) );
  XOR2X1 U202 ( .A(n968), .B(n519), .Y(n1323) );
  XOR2X1 U203 ( .A(n438), .B(n897), .Y(n1245) );
  XOR2X1 U204 ( .A(n1661), .B(n279), .Y(n1399) );
  XOR2X1 U205 ( .A(n1107), .B(n1146), .Y(n718) );
  XOR2X1 U206 ( .A(n311), .B(n1064), .Y(n682) );
  XNOR2X1 U207 ( .A(n979), .B(n980), .Y(n527) );
  XNOR2X1 U208 ( .A(n906), .B(n907), .Y(n446) );
  XOR2X1 U209 ( .A(n1683), .B(n905), .Y(n818) );
  XOR2X1 U210 ( .A(n436), .B(n809), .Y(n887) );
  XOR2X1 U211 ( .A(n357), .B(n735), .Y(n1096) );
  XOR2X1 U212 ( .A(n665), .B(n277), .Y(n1026) );
  XOR2X1 U213 ( .A(n811), .B(n857), .Y(n421) );
  XOR2X1 U214 ( .A(n593), .B(n634), .Y(n501) );
  XOR2X1 U215 ( .A(n359), .B(n1106), .Y(n1165) );
  XOR2X1 U216 ( .A(n737), .B(n775), .Y(n342) );
  XOR2X1 U217 ( .A(n517), .B(n591), .Y(n958) );
  XNOR2X1 U218 ( .A(n1062), .B(n1447), .Y(n685) );
  XOR2X1 U219 ( .A(n631), .B(n1320), .Y(n1004) );
  XOR2X1 U220 ( .A(n667), .B(n702), .Y(n262) );
  XNOR2X1 U221 ( .A(n871), .B(n410), .Y(n1288) );
  XNOR2X1 U222 ( .A(n943), .B(n490), .Y(n1365) );
  XNOR2X1 U223 ( .A(n1080), .B(n329), .Y(n1212) );
  XOR2X1 U224 ( .A(n319), .B(n1391), .Y(n1011) );
  XOR2X1 U225 ( .A(n1662), .B(n643), .Y(n1391) );
  XOR2X1 U226 ( .A(n400), .B(n401), .Y(n399) );
  XNOR2X1 U227 ( .A(n631), .B(n624), .Y(n630) );
  XOR2X1 U228 ( .A(n999), .B(n554), .Y(n613) );
  XNOR2X1 U229 ( .A(n1062), .B(n1063), .Y(n308) );
  XNOR2X1 U230 ( .A(n1136), .B(n1137), .Y(n388) );
  XNOR2X1 U231 ( .A(n966), .B(n1329), .Y(n957) );
  XNOR2X1 U232 ( .A(n1035), .B(n1406), .Y(n1025) );
  XNOR2X1 U233 ( .A(n1212), .B(n1137), .Y(n762) );
  XNOR2X1 U234 ( .A(n895), .B(n1251), .Y(n886) );
  XNOR2X1 U235 ( .A(n1104), .B(n1171), .Y(n1095) );
  XNOR2X1 U236 ( .A(n996), .B(n997), .Y(n552) );
  XOR2X1 U237 ( .A(n1288), .B(n924), .Y(n842) );
  XOR2X1 U238 ( .A(n965), .B(n1329), .Y(n590) );
  XOR2X1 U239 ( .A(n1034), .B(n1406), .Y(n664) );
  XOR2X1 U240 ( .A(n894), .B(n1251), .Y(n808) );
  XOR2X1 U241 ( .A(n1103), .B(n1171), .Y(n734) );
  XNOR2X1 U242 ( .A(n762), .B(n389), .Y(n761) );
  XOR2X1 U243 ( .A(n1034), .B(n1035), .Y(n276) );
  XOR2X1 U244 ( .A(n1103), .B(n1104), .Y(n356) );
  XOR2X1 U245 ( .A(n894), .B(n895), .Y(n435) );
  XOR2X1 U246 ( .A(n1421), .B(n1422), .Y(n1034) );
  XOR2X1 U247 ( .A(n1423), .B(n1424), .Y(n1421) );
  XOR2X1 U248 ( .A(n1047), .B(n1425), .Y(n1424) );
  XOR2X1 U249 ( .A(n1426), .B(n1696), .Y(n1423) );
  XOR2X1 U250 ( .A(n1263), .B(n1264), .Y(n894) );
  XOR2X1 U251 ( .A(n1265), .B(n1266), .Y(n1263) );
  XOR2X1 U252 ( .A(n907), .B(n1267), .Y(n1266) );
  XNOR2X1 U253 ( .A(n1268), .B(n906), .Y(n1265) );
  XOR2X1 U254 ( .A(n1183), .B(n1184), .Y(n1103) );
  XOR2X1 U255 ( .A(n1185), .B(n1186), .Y(n1183) );
  XOR2X1 U256 ( .A(n1187), .B(n1118), .Y(n1186) );
  XNOR2X1 U257 ( .A(n1117), .B(n1188), .Y(n1185) );
  XOR2X1 U258 ( .A(n685), .B(n1055), .Y(n298) );
  XOR2X1 U259 ( .A(n1693), .B(n694), .Y(n1055) );
  XOR2X1 U260 ( .A(n320), .B(n318), .Y(n1070) );
  XOR2X1 U261 ( .A(n808), .B(n809), .Y(n807) );
  XOR2X1 U262 ( .A(n435), .B(n809), .Y(n893) );
  XOR2X1 U263 ( .A(n356), .B(n735), .Y(n1102) );
  XOR2X1 U264 ( .A(n734), .B(n735), .Y(n733) );
  XOR2X1 U265 ( .A(n516), .B(n517), .Y(n515) );
  XOR2X1 U266 ( .A(n590), .B(n517), .Y(n1336) );
  XOR2X1 U267 ( .A(n276), .B(n277), .Y(n275) );
  XOR2X1 U268 ( .A(n664), .B(n277), .Y(n1415) );
  XNOR2X1 U269 ( .A(n624), .B(n625), .Y(n620) );
  XOR2X1 U270 ( .A(n1665), .B(n554), .Y(n625) );
  XOR2X1 U271 ( .A(n664), .B(n665), .Y(n663) );
  XOR2X1 U272 ( .A(n276), .B(n665), .Y(n1033) );
  XOR2X1 U273 ( .A(n1676), .B(n480), .Y(n932) );
  XOR2X1 U274 ( .A(n516), .B(n591), .Y(n964) );
  XOR2X1 U275 ( .A(n590), .B(n591), .Y(n589) );
  XOR2X1 U276 ( .A(n356), .B(n357), .Y(n355) );
  XOR2X1 U277 ( .A(n734), .B(n357), .Y(n1180) );
  XOR2X1 U278 ( .A(n435), .B(n436), .Y(n434) );
  XOR2X1 U279 ( .A(n808), .B(n436), .Y(n1260) );
  XNOR2X1 U280 ( .A(n673), .B(n674), .Y(n672) );
  XOR2X1 U281 ( .A(n468), .B(n457), .Y(n922) );
  XOR2X1 U282 ( .A(n842), .B(n457), .Y(n1296) );
  XNOR2X1 U283 ( .A(n613), .B(n614), .Y(n612) );
  XNOR2X1 U284 ( .A(n287), .B(n288), .Y(n286) );
  XOR2X1 U285 ( .A(n308), .B(n691), .Y(n1061) );
  XNOR2X1 U286 ( .A(n692), .B(n691), .Y(n690) );
  XNOR2X1 U287 ( .A(n623), .B(n622), .Y(n621) );
  XOR2X1 U288 ( .A(n552), .B(n622), .Y(n995) );
  XOR2X1 U289 ( .A(n613), .B(n622), .Y(n1363) );
  XOR2X1 U290 ( .A(n552), .B(n553), .Y(n551) );
  XOR2X1 U291 ( .A(n623), .B(n553), .Y(n1372) );
  XNOR2X1 U292 ( .A(n682), .B(n683), .Y(n681) );
  XOR2X1 U293 ( .A(n388), .B(n389), .Y(n387) );
  XOR2X1 U294 ( .A(n842), .B(n467), .Y(n841) );
  XOR2X1 U295 ( .A(n1116), .B(n366), .Y(n1111) );
  XOR2X1 U296 ( .A(n368), .B(n1119), .Y(n1116) );
  XOR2X1 U297 ( .A(n829), .B(n830), .Y(n828) );
  XOR2X1 U298 ( .A(n831), .B(n456), .Y(n829) );
  XOR2X1 U299 ( .A(n1195), .B(n745), .Y(n1194) );
  XOR2X1 U300 ( .A(n368), .B(n370), .Y(n1195) );
  XOR2X1 U301 ( .A(n1663), .B(n649), .Y(n1397) );
  XOR2X1 U302 ( .A(n1675), .B(n792), .Y(n1242) );
  XOR2X1 U303 ( .A(n1351), .B(n601), .Y(n1350) );
  XOR2X1 U304 ( .A(n529), .B(n528), .Y(n1351) );
  XOR2X1 U305 ( .A(n744), .B(n367), .Y(n1112) );
  XOR2X1 U306 ( .A(n1275), .B(n817), .Y(n1274) );
  XOR2X1 U307 ( .A(n448), .B(n449), .Y(n1275) );
  XOR2X1 U308 ( .A(n1699), .B(n718), .Y(n1162) );
  XOR2X1 U309 ( .A(n1043), .B(n674), .Y(n1042) );
  XOR2X1 U310 ( .A(n298), .B(n299), .Y(n297) );
  XOR2X1 U311 ( .A(n1287), .B(n916), .Y(n1286) );
  XOR2X1 U312 ( .A(n831), .B(n830), .Y(n1287) );
  XOR2X1 U313 ( .A(n539), .B(n540), .Y(n538) );
  XNOR2X1 U314 ( .A(n541), .B(n542), .Y(n539) );
  XOR2X1 U315 ( .A(n1690), .B(n709), .Y(n708) );
  XOR2X1 U316 ( .A(n1677), .B(n783), .Y(n782) );
  XNOR2X1 U317 ( .A(n401), .B(n709), .Y(n1078) );
  XOR2X1 U318 ( .A(n479), .B(n783), .Y(n869) );
  XOR2X1 U319 ( .A(n988), .B(n614), .Y(n987) );
  XNOR2X1 U320 ( .A(n541), .B(n540), .Y(n988) );
  XNOR2X1 U321 ( .A(n320), .B(n321), .Y(n316) );
  XNOR2X1 U322 ( .A(n448), .B(n449), .Y(n444) );
  XOR2X1 U323 ( .A(n1669), .B(n566), .Y(n565) );
  XNOR2X1 U324 ( .A(n411), .B(n410), .Y(n406) );
  XNOR2X1 U325 ( .A(n491), .B(n490), .Y(n486) );
  XNOR2X1 U326 ( .A(n330), .B(n329), .Y(n325) );
  XOR2X1 U327 ( .A(n448), .B(n447), .Y(n815) );
  XOR2X1 U328 ( .A(n1676), .B(n481), .Y(n477) );
  XOR2X1 U329 ( .A(n884), .B(n885), .Y(n426) );
  XOR2X1 U330 ( .A(n886), .B(n887), .Y(n884) );
  XOR2X1 U331 ( .A(n1352), .B(n1340), .Y(n529) );
  XOR2X1 U332 ( .A(n1355), .B(n1356), .Y(n1352) );
  XNOR2X1 U333 ( .A(n999), .B(n557), .Y(n1355) );
  XNOR2X1 U334 ( .A(n554), .B(n624), .Y(n1356) );
  XOR2X1 U335 ( .A(n529), .B(n530), .Y(n525) );
  XNOR2X1 U336 ( .A(n531), .B(n532), .Y(n530) );
  XOR2X1 U337 ( .A(n368), .B(n369), .Y(n364) );
  XNOR2X1 U338 ( .A(n370), .B(n371), .Y(n369) );
  XOR2X1 U339 ( .A(n656), .B(n1663), .Y(n655) );
  XOR2X1 U340 ( .A(n259), .B(n1663), .Y(n1017) );
  XOR2X1 U341 ( .A(n800), .B(n1675), .Y(n799) );
  XOR2X1 U342 ( .A(n726), .B(n1699), .Y(n725) );
  XOR2X1 U343 ( .A(n583), .B(n1668), .Y(n582) );
  XOR2X1 U344 ( .A(n754), .B(n1688), .Y(n1208) );
  XNOR2X1 U345 ( .A(n566), .B(n941), .Y(n940) );
  XNOR2X1 U346 ( .A(n298), .B(n1054), .Y(n1053) );
  XOR2X1 U347 ( .A(n3), .B(n744), .Y(n742) );
  XNOR2X1 U348 ( .A(n368), .B(n745), .Y(n3) );
  XOR2X1 U349 ( .A(n289), .B(n290), .Y(n285) );
  XOR2X1 U350 ( .A(n1659), .B(n291), .Y(n290) );
  XOR2X1 U351 ( .A(n499), .B(n500), .Y(n495) );
  XOR2X1 U352 ( .A(n1671), .B(n501), .Y(n500) );
  XOR2X1 U353 ( .A(n419), .B(n420), .Y(n415) );
  XOR2X1 U354 ( .A(n1682), .B(n421), .Y(n420) );
  XOR2X1 U355 ( .A(n1339), .B(n1340), .Y(n965) );
  XOR2X1 U356 ( .A(n1341), .B(n1342), .Y(n1339) );
  XOR2X1 U357 ( .A(n1343), .B(n980), .Y(n1342) );
  XOR2X1 U358 ( .A(n979), .B(n1697), .Y(n1341) );
  INVX1 U359 ( .A(n956), .Y(n1669) );
  INVX1 U360 ( .A(n1094), .Y(n1690) );
  INVX1 U361 ( .A(n1024), .Y(n1656) );
  INVX1 U362 ( .A(n885), .Y(n1677) );
  INVX1 U363 ( .A(n1405), .Y(n1661) );
  INVX1 U364 ( .A(n469), .Y(n1684) );
  INVX1 U365 ( .A(n1440), .Y(n1693) );
  INVX1 U366 ( .A(n933), .Y(n1676) );
  INVX1 U367 ( .A(n1344), .Y(n1697) );
  INVX1 U368 ( .A(n1046), .Y(n1696) );
  XNOR2X1 U369 ( .A(n1288), .B(n923), .Y(n831) );
  XNOR2X1 U370 ( .A(n468), .B(n467), .Y(n466) );
  XNOR2X1 U371 ( .A(n248), .B(n249), .Y(n247) );
  XOR2X1 U372 ( .A(n969), .B(n1320), .Y(n575) );
  XNOR2X1 U373 ( .A(n1268), .B(n1267), .Y(n817) );
  XNOR2X1 U374 ( .A(n1117), .B(n1118), .Y(n366) );
  XOR2X1 U375 ( .A(n1200), .B(n379), .Y(n1135) );
  XOR2X1 U376 ( .A(n327), .B(n328), .Y(n326) );
  XOR2X1 U377 ( .A(n1672), .B(n977), .Y(n602) );
  XOR2X1 U378 ( .A(n1384), .B(n941), .Y(n1473) );
  XOR2X1 U379 ( .A(n479), .B(n885), .Y(n1235) );
  XNOR2X1 U380 ( .A(n1426), .B(n1425), .Y(n673) );
  XOR2X1 U381 ( .A(n488), .B(n489), .Y(n487) );
  XOR2X1 U382 ( .A(n408), .B(n409), .Y(n407) );
  XNOR2X1 U383 ( .A(n318), .B(n319), .Y(n317) );
  XOR2X1 U384 ( .A(n479), .B(n480), .Y(n478) );
  XOR2X1 U385 ( .A(n456), .B(n457), .Y(n455) );
  XOR2X1 U386 ( .A(n1054), .B(n691), .Y(n1445) );
  XOR2X1 U387 ( .A(n378), .B(n389), .Y(n1124) );
  XOR2X1 U388 ( .A(n446), .B(n447), .Y(n445) );
  XOR2X1 U389 ( .A(n378), .B(n379), .Y(n377) );
  XOR2X1 U390 ( .A(n1668), .B(n575), .Y(n1319) );
  XOR2X1 U391 ( .A(n527), .B(n528), .Y(n526) );
  XOR2X1 U392 ( .A(n366), .B(n367), .Y(n365) );
  XOR2X1 U393 ( .A(n1144), .B(n398), .Y(n1143) );
  XOR2X1 U394 ( .A(n467), .B(n916), .Y(n915) );
  XOR2X1 U395 ( .A(n1043), .B(n673), .Y(n1433) );
  XOR2X1 U396 ( .A(n328), .B(n1080), .Y(n1077) );
  XOR2X1 U397 ( .A(n489), .B(n943), .Y(n939) );
  XNOR2X1 U398 ( .A(n279), .B(n666), .Y(n662) );
  XOR2X1 U399 ( .A(n667), .B(n1664), .Y(n666) );
  XNOR2X1 U400 ( .A(n438), .B(n810), .Y(n806) );
  XOR2X1 U401 ( .A(n811), .B(n1678), .Y(n810) );
  XNOR2X1 U402 ( .A(n897), .B(n1269), .Y(n1259) );
  XOR2X1 U403 ( .A(n811), .B(n1686), .Y(n1269) );
  XNOR2X1 U404 ( .A(n359), .B(n736), .Y(n732) );
  XOR2X1 U405 ( .A(n737), .B(n1700), .Y(n736) );
  XNOR2X1 U406 ( .A(n1106), .B(n1189), .Y(n1179) );
  XOR2X1 U407 ( .A(n737), .B(n1692), .Y(n1189) );
  XOR2X1 U408 ( .A(n409), .B(n871), .Y(n868) );
  XOR2X1 U409 ( .A(n941), .B(n1669), .Y(n1313) );
  XOR2X1 U410 ( .A(n401), .B(n1690), .Y(n1155) );
  XOR2X1 U411 ( .A(n1405), .B(n1428), .Y(n1414) );
  XOR2X1 U412 ( .A(n667), .B(n1658), .Y(n1428) );
  INVX1 U413 ( .A(n1037), .Y(n1657) );
  INVX1 U414 ( .A(n898), .Y(n1679) );
  INVX1 U415 ( .A(n1107), .Y(n1691) );
  INVX1 U416 ( .A(n969), .Y(n1670) );
  BUFX2 U417 ( .A(n244), .Y(n97) );
  BUFX2 U418 ( .A(n244), .Y(n88) );
  BUFX2 U419 ( .A(n244), .Y(n85) );
  BUFX2 U420 ( .A(n244), .Y(n91) );
  BUFX2 U421 ( .A(n244), .Y(n96) );
  BUFX2 U422 ( .A(n242), .Y(n101) );
  BUFX2 U423 ( .A(n147), .Y(n108) );
  BUFX2 U424 ( .A(n107), .Y(n147) );
  BUFX2 U425 ( .A(n242), .Y(n107) );
  INVX1 U426 ( .A(n1485), .Y(n1703) );
  AOI21X1 U427 ( .A0(n1476), .A1(n1477), .B0(n1489), .Y(n1474) );
  NAND2X1 U428 ( .A(n1148), .B(n860), .Y(n205) );
  NAND2X1 U429 ( .A(n862), .B(n860), .Y(n204) );
  NAND2X1 U430 ( .A(n1469), .B(n860), .Y(n201) );
  INVX1 U431 ( .A(n1475), .Y(n1704) );
  INVX1 U432 ( .A(n1476), .Y(n1707) );
  BUFX2 U433 ( .A(n202), .Y(n1634) );
  INVX1 U434 ( .A(n1477), .Y(n1705) );
  BUFX2 U435 ( .A(n202), .Y(n1635) );
  BUFX2 U436 ( .A(n202), .Y(n1636) );
  XOR2X1 U437 ( .A(n261), .B(n268), .Y(n249) );
  XOR2X1 U438 ( .A(n348), .B(n341), .Y(n328) );
  XOR2X1 U439 ( .A(n877), .B(n418), .Y(n885) );
  XOR2X1 U440 ( .A(n949), .B(n497), .Y(n956) );
  XOR2X1 U441 ( .A(n1086), .B(n337), .Y(n1094) );
  XNOR2X1 U442 ( .A(n314), .B(n243), .Y(n1440) );
  XNOR2X1 U443 ( .A(n1028), .B(n1658), .Y(n1037) );
  XNOR2X1 U444 ( .A(n970), .B(n1686), .Y(n898) );
  XNOR2X1 U445 ( .A(n1163), .B(n1692), .Y(n1107) );
  XOR2X1 U446 ( .A(n510), .B(n594), .Y(n969) );
  XNOR2X1 U447 ( .A(n543), .B(n569), .Y(n1344) );
  XNOR2X1 U448 ( .A(n523), .B(n484), .Y(n1405) );
  XOR2X1 U449 ( .A(n1427), .B(n251), .Y(n1046) );
  XNOR2X1 U450 ( .A(n427), .B(n1244), .Y(n409) );
  XNOR2X1 U451 ( .A(n507), .B(n1322), .Y(n489) );
  XOR2X1 U452 ( .A(n1140), .B(n1685), .Y(n469) );
  XOR2X1 U453 ( .A(n1437), .B(n258), .Y(n1024) );
  XNOR2X1 U454 ( .A(n1114), .B(n1115), .Y(n744) );
  XNOR2X1 U455 ( .A(n1140), .B(n855), .Y(n933) );
  XNOR2X1 U456 ( .A(n788), .B(n942), .Y(n491) );
  XNOR2X1 U457 ( .A(n879), .B(n870), .Y(n411) );
  XNOR2X1 U458 ( .A(n1088), .B(n1079), .Y(n330) );
  XNOR2X1 U459 ( .A(n697), .B(n637), .Y(n624) );
  XOR2X1 U460 ( .A(n475), .B(n404), .Y(n694) );
  XOR2X1 U461 ( .A(n1201), .B(n777), .Y(n764) );
  XOR2X1 U462 ( .A(n854), .B(n1681), .Y(n472) );
  XOR2X1 U463 ( .A(n853), .B(n859), .Y(n844) );
  XOR2X1 U464 ( .A(n633), .B(n567), .Y(n557) );
  XOR2X1 U465 ( .A(n852), .B(n935), .Y(n926) );
  XOR2X1 U466 ( .A(n774), .B(n710), .Y(n390) );
  XOR2X1 U467 ( .A(n1071), .B(n484), .Y(n1064) );
  XNOR2X1 U468 ( .A(n641), .B(n251), .Y(n318) );
  XOR2X1 U469 ( .A(n1695), .B(n562), .Y(n554) );
  XNOR2X1 U470 ( .A(n545), .B(n1358), .Y(n982) );
  XOR2X1 U471 ( .A(n821), .B(n859), .Y(n809) );
  XOR2X1 U472 ( .A(n747), .B(n777), .Y(n735) );
  XNOR2X1 U473 ( .A(n978), .B(n567), .Y(n517) );
  XOR2X1 U474 ( .A(n283), .B(n243), .Y(n277) );
  XOR2X1 U475 ( .A(n1674), .B(n785), .Y(n857) );
  XOR2X1 U476 ( .A(n1667), .B(n569), .Y(n634) );
  XOR2X1 U477 ( .A(n442), .B(n404), .Y(n665) );
  XOR2X1 U478 ( .A(n417), .B(n879), .Y(n480) );
  XOR2X1 U479 ( .A(n825), .B(n567), .Y(n532) );
  XOR2X1 U480 ( .A(n604), .B(n637), .Y(n591) );
  XOR2X1 U481 ( .A(n1698), .B(n712), .Y(n775) );
  XNOR2X1 U482 ( .A(n756), .B(n1203), .Y(n1119) );
  XOR2X1 U483 ( .A(n1114), .B(n710), .Y(n357) );
  XOR2X1 U484 ( .A(n1048), .B(n1236), .Y(n436) );
  XOR2X1 U485 ( .A(n280), .B(n270), .Y(n667) );
  XOR2X1 U486 ( .A(n439), .B(n429), .Y(n811) );
  XOR2X1 U487 ( .A(n360), .B(n350), .Y(n737) );
  XOR2X1 U488 ( .A(n520), .B(n509), .Y(n593) );
  XOR2X1 U489 ( .A(n935), .B(n859), .Y(n408) );
  XOR2X1 U490 ( .A(n498), .B(n788), .Y(n1320) );
  XOR2X1 U491 ( .A(n396), .B(n1655), .Y(n311) );
  XOR2X1 U492 ( .A(n597), .B(n562), .Y(n519) );
  XOR2X1 U493 ( .A(n1147), .B(n1689), .Y(n393) );
  XOR2X1 U494 ( .A(n833), .B(n935), .Y(n909) );
  XOR2X1 U495 ( .A(n822), .B(n935), .Y(n897) );
  XOR2X1 U496 ( .A(n768), .B(n1666), .Y(n999) );
  XOR2X1 U497 ( .A(n1662), .B(n333), .Y(n702) );
  XNOR2X1 U498 ( .A(n463), .B(n641), .Y(n1047) );
  XNOR2X1 U499 ( .A(n556), .B(n577), .Y(n1343) );
  XOR2X1 U500 ( .A(n452), .B(n404), .Y(n1044) );
  XOR2X1 U501 ( .A(n381), .B(n777), .Y(n1115) );
  XOR2X1 U502 ( .A(n471), .B(n785), .Y(n1267) );
  XOR2X1 U503 ( .A(n1685), .B(n785), .Y(n410) );
  XOR2X1 U504 ( .A(n562), .B(n569), .Y(n490) );
  XOR2X1 U505 ( .A(n535), .B(n484), .Y(n1418) );
  XOR2X1 U506 ( .A(n1689), .B(n712), .Y(n329) );
  XOR2X1 U507 ( .A(n1203), .B(n720), .Y(n1080) );
  XNOR2X1 U508 ( .A(n372), .B(n1655), .Y(n279) );
  XNOR2X1 U509 ( .A(n459), .B(n858), .Y(n820) );
  XOR2X1 U510 ( .A(n1358), .B(n577), .Y(n943) );
  XNOR2X1 U511 ( .A(n834), .B(n417), .Y(n906) );
  XOR2X1 U512 ( .A(n832), .B(n859), .Y(n905) );
  XOR2X1 U513 ( .A(n1125), .B(n720), .Y(n1188) );
  XOR2X1 U514 ( .A(n755), .B(n338), .Y(n1118) );
  XOR2X1 U515 ( .A(n1126), .B(n1689), .Y(n371) );
  XOR2X1 U516 ( .A(n294), .B(n243), .Y(n1409) );
  XOR2X1 U517 ( .A(n1128), .B(n710), .Y(n1174) );
  XOR2X1 U518 ( .A(n392), .B(n712), .Y(n1187) );
  XNOR2X1 U519 ( .A(n300), .B(n333), .Y(n1426) );
  XOR2X1 U520 ( .A(n748), .B(n1694), .Y(n1106) );
  XOR2X1 U521 ( .A(n546), .B(n788), .Y(n980) );
  XOR2X1 U522 ( .A(n616), .B(n637), .Y(n977) );
  XOR2X1 U523 ( .A(n845), .B(n879), .Y(n907) );
  XNOR2X1 U524 ( .A(n302), .B(n1419), .Y(n676) );
  XOR2X1 U525 ( .A(n609), .B(n562), .Y(n606) );
  XOR2X1 U526 ( .A(n1201), .B(n1144), .Y(n400) );
  XOR2X1 U527 ( .A(n1071), .B(n1072), .Y(n320) );
  XOR2X1 U528 ( .A(n765), .B(n1088), .Y(n1117) );
  XOR2X1 U529 ( .A(n773), .B(n1694), .Y(n1200) );
  XOR2X1 U530 ( .A(n1448), .B(n1449), .Y(n1062) );
  XOR2X1 U531 ( .A(n641), .B(n404), .Y(n1448) );
  XOR2X1 U532 ( .A(n243), .B(n251), .Y(n1449) );
  XOR2X1 U533 ( .A(n989), .B(n498), .Y(n979) );
  XOR2X1 U534 ( .A(n910), .B(n1685), .Y(n438) );
  XOR2X1 U535 ( .A(n605), .B(n1666), .Y(n968) );
  XOR2X1 U536 ( .A(n1113), .B(n1689), .Y(n359) );
  XOR2X1 U537 ( .A(n1682), .B(n427), .Y(n1277) );
  XOR2X1 U538 ( .A(n1671), .B(n507), .Y(n1353) );
  XNOR2X1 U539 ( .A(n1455), .B(n1456), .Y(n1063) );
  XOR2X1 U540 ( .A(n1458), .B(n1459), .Y(n1455) );
  XOR2X1 U541 ( .A(n1457), .B(n249), .Y(n1456) );
  XOR2X1 U542 ( .A(n1437), .B(n1660), .Y(n1458) );
  XOR2X1 U543 ( .A(n1289), .B(n1290), .Y(n923) );
  XOR2X1 U544 ( .A(n1236), .B(n417), .Y(n1289) );
  XOR2X1 U545 ( .A(n879), .B(n859), .Y(n1290) );
  XOR2X1 U546 ( .A(n1213), .B(n1214), .Y(n1136) );
  XNOR2X1 U547 ( .A(n338), .B(n710), .Y(n1213) );
  XOR2X1 U548 ( .A(n1088), .B(n777), .Y(n1214) );
  XOR2X1 U549 ( .A(n442), .B(n1409), .Y(n291) );
  XNOR2X1 U550 ( .A(n1297), .B(n1298), .Y(n924) );
  XOR2X1 U551 ( .A(n1300), .B(n1301), .Y(n1297) );
  XOR2X1 U552 ( .A(n1299), .B(n1277), .Y(n1298) );
  XOR2X1 U553 ( .A(n1674), .B(n418), .Y(n1301) );
  XNOR2X1 U554 ( .A(n1220), .B(n1221), .Y(n1137) );
  XOR2X1 U555 ( .A(n1094), .B(n1223), .Y(n1220) );
  XOR2X1 U556 ( .A(n1222), .B(n328), .Y(n1221) );
  XOR2X1 U557 ( .A(n1698), .B(n338), .Y(n1223) );
  XOR2X1 U558 ( .A(n283), .B(n1044), .Y(n674) );
  XNOR2X1 U559 ( .A(n1337), .B(n1338), .Y(n1329) );
  XOR2X1 U560 ( .A(n577), .B(n569), .Y(n1337) );
  XOR2X1 U561 ( .A(n606), .B(n982), .Y(n1338) );
  XOR2X1 U562 ( .A(n333), .B(n251), .Y(n1457) );
  XOR2X1 U563 ( .A(n250), .B(n251), .Y(n246) );
  XOR2X1 U564 ( .A(n252), .B(n1655), .Y(n250) );
  XNOR2X1 U565 ( .A(n1416), .B(n1417), .Y(n1406) );
  XOR2X1 U566 ( .A(n1420), .B(n333), .Y(n1416) );
  XOR2X1 U567 ( .A(n676), .B(n1418), .Y(n1417) );
  XNOR2X1 U568 ( .A(n1261), .B(n1262), .Y(n1251) );
  XOR2X1 U569 ( .A(n794), .B(n785), .Y(n1261) );
  XOR2X1 U570 ( .A(n909), .B(n820), .Y(n1262) );
  XNOR2X1 U571 ( .A(n1181), .B(n1182), .Y(n1171) );
  XOR2X1 U572 ( .A(n720), .B(n712), .Y(n1181) );
  XOR2X1 U573 ( .A(n1119), .B(n371), .Y(n1182) );
  XOR2X1 U574 ( .A(n338), .B(n1079), .Y(n709) );
  XOR2X1 U575 ( .A(n417), .B(n870), .Y(n783) );
  XOR2X1 U576 ( .A(n419), .B(n877), .Y(n876) );
  XOR2X1 U577 ( .A(n1460), .B(n1461), .Y(n1447) );
  XOR2X1 U578 ( .A(n1420), .B(n484), .Y(n1460) );
  XOR2X1 U579 ( .A(n1655), .B(n333), .Y(n1461) );
  XOR2X1 U580 ( .A(n910), .B(n1254), .Y(n449) );
  XOR2X1 U581 ( .A(n879), .B(n785), .Y(n1299) );
  XOR2X1 U582 ( .A(n1088), .B(n712), .Y(n1222) );
  XOR2X1 U583 ( .A(n1667), .B(n498), .Y(n1376) );
  XNOR2X1 U584 ( .A(n1407), .B(n1408), .Y(n1035) );
  XOR2X1 U585 ( .A(n641), .B(n251), .Y(n1407) );
  XOR2X1 U586 ( .A(n1409), .B(n1044), .Y(n1408) );
  XOR2X1 U587 ( .A(n747), .B(n1174), .Y(n370) );
  XNOR2X1 U588 ( .A(n1172), .B(n1173), .Y(n1104) );
  XNOR2X1 U589 ( .A(n338), .B(n1088), .Y(n1172) );
  XOR2X1 U590 ( .A(n1174), .B(n1115), .Y(n1173) );
  XNOR2X1 U591 ( .A(n768), .B(n1385), .Y(n631) );
  XOR2X1 U592 ( .A(n605), .B(n606), .Y(n531) );
  XOR2X1 U593 ( .A(n339), .B(n1086), .Y(n1085) );
  XNOR2X1 U594 ( .A(n1252), .B(n1253), .Y(n895) );
  XNOR2X1 U595 ( .A(n417), .B(n879), .Y(n1252) );
  XOR2X1 U596 ( .A(n905), .B(n1254), .Y(n1253) );
  XOR2X1 U597 ( .A(n249), .B(n1436), .Y(n1422) );
  XOR2X1 U598 ( .A(n258), .B(n1663), .Y(n1436) );
  XOR2X1 U599 ( .A(n1277), .B(n1278), .Y(n1264) );
  XOR2X1 U600 ( .A(n418), .B(n1675), .Y(n1278) );
  XOR2X1 U601 ( .A(n1353), .B(n1354), .Y(n1340) );
  XOR2X1 U602 ( .A(n497), .B(n1668), .Y(n1354) );
  XOR2X1 U603 ( .A(n328), .B(n1197), .Y(n1184) );
  XOR2X1 U604 ( .A(n337), .B(n1699), .Y(n1197) );
  XOR2X1 U605 ( .A(n499), .B(n949), .Y(n948) );
  XOR2X1 U606 ( .A(n800), .B(n418), .Y(n1250) );
  XOR2X1 U607 ( .A(n877), .B(n417), .Y(n1300) );
  XOR2X1 U608 ( .A(n498), .B(n942), .Y(n566) );
  XNOR2X1 U609 ( .A(n333), .B(n643), .Y(n252) );
  XOR2X1 U610 ( .A(n1662), .B(n258), .Y(n1459) );
  XOR2X1 U611 ( .A(n656), .B(n258), .Y(n1404) );
  XOR2X1 U612 ( .A(n836), .B(n1681), .Y(n1254) );
  XOR2X1 U613 ( .A(n1366), .B(n1367), .Y(n996) );
  XNOR2X1 U614 ( .A(n637), .B(n788), .Y(n1366) );
  XOR2X1 U615 ( .A(n567), .B(n498), .Y(n1367) );
  XOR2X1 U616 ( .A(n310), .B(n1662), .Y(n1425) );
  XOR2X1 U617 ( .A(n1314), .B(n1667), .Y(n1312) );
  XOR2X1 U618 ( .A(n491), .B(n637), .Y(n1314) );
  XOR2X1 U619 ( .A(n583), .B(n497), .Y(n1328) );
  XOR2X1 U620 ( .A(n726), .B(n337), .Y(n1170) );
  XOR2X1 U621 ( .A(n935), .B(n1674), .Y(n871) );
  XOR2X1 U622 ( .A(n754), .B(n755), .Y(n753) );
  XOR2X1 U623 ( .A(n925), .B(n926), .Y(n921) );
  XOR2X1 U624 ( .A(n927), .B(n844), .Y(n925) );
  XOR2X1 U625 ( .A(n933), .B(n853), .Y(n1307) );
  XOR2X1 U626 ( .A(n632), .B(n633), .Y(n629) );
  XNOR2X1 U627 ( .A(n562), .B(n634), .Y(n632) );
  XOR2X1 U628 ( .A(n927), .B(n1674), .Y(n1268) );
  XOR2X1 U629 ( .A(n1386), .B(n567), .Y(n1381) );
  XOR2X1 U630 ( .A(n1358), .B(n634), .Y(n1386) );
  XOR2X1 U631 ( .A(n615), .B(n553), .Y(n611) );
  XNOR2X1 U632 ( .A(n541), .B(n616), .Y(n615) );
  XOR2X1 U633 ( .A(n1687), .B(n380), .Y(n376) );
  XOR2X1 U634 ( .A(n381), .B(n382), .Y(n380) );
  XOR2X1 U635 ( .A(n1687), .B(n1127), .Y(n1123) );
  XOR2X1 U636 ( .A(n1128), .B(n382), .Y(n1127) );
  XOR2X1 U637 ( .A(n258), .B(n649), .Y(n648) );
  XOR2X1 U638 ( .A(n642), .B(n248), .Y(n639) );
  XOR2X1 U639 ( .A(n252), .B(n243), .Y(n642) );
  XOR2X1 U640 ( .A(n418), .B(n792), .Y(n791) );
  XOR2X1 U641 ( .A(n851), .B(n481), .Y(n850) );
  XNOR2X1 U642 ( .A(n854), .B(n855), .Y(n851) );
  XOR2X1 U643 ( .A(n337), .B(n718), .Y(n717) );
  XOR2X1 U644 ( .A(n1383), .B(n1384), .Y(n1382) );
  XNOR2X1 U645 ( .A(n633), .B(n1385), .Y(n1383) );
  XOR2X1 U646 ( .A(n400), .B(n772), .Y(n771) );
  XOR2X1 U647 ( .A(n773), .B(n774), .Y(n772) );
  XOR2X1 U648 ( .A(n400), .B(n1229), .Y(n1228) );
  XOR2X1 U649 ( .A(n1147), .B(n774), .Y(n1229) );
  XOR2X1 U650 ( .A(n320), .B(n701), .Y(n700) );
  XOR2X1 U651 ( .A(n475), .B(n314), .Y(n701) );
  XOR2X1 U652 ( .A(n339), .B(n1164), .Y(n1161) );
  XNOR2X1 U653 ( .A(n341), .B(n712), .Y(n1164) );
  XOR2X1 U654 ( .A(n1209), .B(n1210), .Y(n754) );
  XOR2X1 U655 ( .A(n393), .B(n1211), .Y(n1210) );
  XOR2X1 U656 ( .A(n1129), .B(n1200), .Y(n1209) );
  XOR2X1 U657 ( .A(n1128), .B(n381), .Y(n1211) );
  XOR2X1 U658 ( .A(n1072), .B(n1467), .Y(n1466) );
  XOR2X1 U659 ( .A(n314), .B(n321), .Y(n1467) );
  XOR2X1 U660 ( .A(n1045), .B(n287), .Y(n1041) );
  XOR2X1 U661 ( .A(n289), .B(n523), .Y(n1045) );
  XOR2X1 U662 ( .A(n419), .B(n1243), .Y(n1241) );
  XOR2X1 U663 ( .A(n1244), .B(n785), .Y(n1243) );
  XOR2X1 U664 ( .A(n1446), .B(n682), .Y(n1444) );
  XOR2X1 U665 ( .A(n685), .B(n452), .Y(n1446) );
  XOR2X1 U666 ( .A(n499), .B(n1321), .Y(n1318) );
  XOR2X1 U667 ( .A(n1322), .B(n569), .Y(n1321) );
  XOR2X1 U668 ( .A(n684), .B(n299), .Y(n680) );
  XOR2X1 U669 ( .A(n685), .B(n294), .Y(n684) );
  XOR2X1 U670 ( .A(n1660), .B(n1012), .Y(n1010) );
  XOR2X1 U671 ( .A(n484), .B(n249), .Y(n1012) );
  XOR2X1 U672 ( .A(n675), .B(n288), .Y(n671) );
  XOR2X1 U673 ( .A(n289), .B(n442), .Y(n675) );
  XNOR2X1 U674 ( .A(n1373), .B(n1374), .Y(n997) );
  XOR2X1 U675 ( .A(n1375), .B(n1353), .Y(n1374) );
  XOR2X1 U676 ( .A(n956), .B(n1376), .Y(n1373) );
  XOR2X1 U677 ( .A(n788), .B(n569), .Y(n1375) );
  XOR2X1 U678 ( .A(n419), .B(n793), .Y(n790) );
  XOR2X1 U679 ( .A(n794), .B(n427), .Y(n793) );
  XOR2X1 U680 ( .A(n1064), .B(n1065), .Y(n1060) );
  XOR2X1 U681 ( .A(n300), .B(n694), .Y(n1065) );
  XOR2X1 U682 ( .A(n311), .B(n693), .Y(n689) );
  XOR2X1 U683 ( .A(n463), .B(n694), .Y(n693) );
  XOR2X1 U684 ( .A(n499), .B(n576), .Y(n573) );
  XOR2X1 U685 ( .A(n577), .B(n507), .Y(n576) );
  XOR2X1 U686 ( .A(n501), .B(n950), .Y(n947) );
  XOR2X1 U687 ( .A(n788), .B(n507), .Y(n950) );
  XOR2X1 U688 ( .A(n339), .B(n719), .Y(n716) );
  XOR2X1 U689 ( .A(n720), .B(n348), .Y(n719) );
  XOR2X1 U690 ( .A(n259), .B(n1398), .Y(n1396) );
  XOR2X1 U691 ( .A(n333), .B(n261), .Y(n1398) );
  XOR2X1 U692 ( .A(n1681), .B(n784), .Y(n781) );
  XOR2X1 U693 ( .A(n785), .B(n408), .Y(n784) );
  XOR2X1 U694 ( .A(n1673), .B(n458), .Y(n454) );
  XOR2X1 U695 ( .A(n459), .B(n460), .Y(n458) );
  XOR2X1 U696 ( .A(n1673), .B(n917), .Y(n914) );
  XOR2X1 U697 ( .A(n833), .B(n460), .Y(n917) );
  XOR2X1 U698 ( .A(n289), .B(n1434), .Y(n1432) );
  XOR2X1 U699 ( .A(n283), .B(n291), .Y(n1434) );
  XOR2X1 U700 ( .A(n541), .B(n1364), .Y(n1362) );
  XOR2X1 U701 ( .A(n825), .B(n542), .Y(n1364) );
  XOR2X1 U702 ( .A(n339), .B(n340), .Y(n335) );
  XOR2X1 U703 ( .A(n341), .B(n342), .Y(n340) );
  XOR2X1 U704 ( .A(n259), .B(n260), .Y(n256) );
  XOR2X1 U705 ( .A(n261), .B(n262), .Y(n260) );
  XOR2X1 U706 ( .A(n529), .B(n603), .Y(n599) );
  XOR2X1 U707 ( .A(n604), .B(n531), .Y(n603) );
  XOR2X1 U708 ( .A(n259), .B(n650), .Y(n647) );
  XOR2X1 U709 ( .A(n268), .B(n1662), .Y(n650) );
  XOR2X1 U710 ( .A(n1237), .B(n1674), .Y(n1234) );
  XOR2X1 U711 ( .A(n411), .B(n859), .Y(n1237) );
  XOR2X1 U712 ( .A(n1157), .B(n1698), .Y(n1154) );
  XOR2X1 U713 ( .A(n330), .B(n777), .Y(n1157) );
  INVX1 U714 ( .A(n641), .Y(n1660) );
  INVX1 U715 ( .A(n1419), .Y(n1655) );
  INVX1 U716 ( .A(n794), .Y(n1674) );
  INVX1 U717 ( .A(n720), .Y(n1698) );
  INVX1 U718 ( .A(n1420), .Y(n1662) );
  INVX1 U719 ( .A(n577), .Y(n1667) );
  INVX1 U720 ( .A(n858), .Y(n1685) );
  INVX1 U721 ( .A(n1358), .Y(n1666) );
  INVX1 U722 ( .A(n1203), .Y(n1694) );
  INVX1 U723 ( .A(n1437), .Y(n1663) );
  INVX1 U724 ( .A(n1156), .Y(n1689) );
  INVX1 U725 ( .A(n877), .Y(n1675) );
  INVX1 U726 ( .A(n1236), .Y(n1681) );
  INVX1 U727 ( .A(n1086), .Y(n1699) );
  INVX1 U728 ( .A(n949), .Y(n1668) );
  INVX1 U729 ( .A(n1322), .Y(n1671) );
  INVX1 U730 ( .A(n1244), .Y(n1682) );
  INVX1 U731 ( .A(n658), .Y(n1658) );
  INVX1 U732 ( .A(n802), .Y(n1686) );
  INVX1 U733 ( .A(n728), .Y(n1692) );
  INVX1 U734 ( .A(n1005), .Y(n1695) );
  XNOR2X1 U735 ( .A(n562), .B(n567), .Y(n941) );
  XOR2X1 U736 ( .A(n1156), .B(n710), .Y(n401) );
  XNOR2X1 U737 ( .A(n294), .B(n302), .Y(n1054) );
  XOR2X1 U738 ( .A(n1694), .B(n777), .Y(n327) );
  XOR2X1 U739 ( .A(n484), .B(n404), .Y(n248) );
  XOR2X1 U740 ( .A(n471), .B(n845), .Y(n457) );
  XOR2X1 U741 ( .A(n1701), .B(n310), .Y(n691) );
  XOR2X1 U742 ( .A(n546), .B(n556), .Y(n622) );
  XOR2X1 U743 ( .A(n1665), .B(n543), .Y(n553) );
  XOR2X1 U744 ( .A(n1125), .B(n755), .Y(n389) );
  XOR2X1 U745 ( .A(n1680), .B(n834), .Y(n467) );
  XOR2X1 U746 ( .A(n338), .B(n1088), .Y(n1146) );
  XOR2X1 U747 ( .A(n1655), .B(n243), .Y(n319) );
  XNOR2X1 U748 ( .A(n819), .B(n820), .Y(n447) );
  XNOR2X1 U749 ( .A(n821), .B(n822), .Y(n819) );
  XNOR2X1 U750 ( .A(n1236), .B(n1685), .Y(n479) );
  XOR2X1 U751 ( .A(n637), .B(n1666), .Y(n488) );
  XOR2X1 U752 ( .A(n1688), .B(n392), .Y(n379) );
  XNOR2X1 U753 ( .A(n337), .B(n338), .Y(n336) );
  XOR2X1 U754 ( .A(n702), .B(n703), .Y(n699) );
  XOR2X1 U755 ( .A(n1655), .B(n404), .Y(n703) );
  XOR2X1 U756 ( .A(n852), .B(n853), .Y(n481) );
  XOR2X1 U757 ( .A(n604), .B(n597), .Y(n528) );
  XOR2X1 U758 ( .A(n1113), .B(n748), .Y(n367) );
  XNOR2X1 U759 ( .A(n497), .B(n498), .Y(n496) );
  XNOR2X1 U760 ( .A(n1145), .B(n1146), .Y(n398) );
  XNOR2X1 U761 ( .A(n773), .B(n1147), .Y(n1145) );
  XOR2X1 U762 ( .A(n452), .B(n535), .Y(n299) );
  XOR2X1 U763 ( .A(n836), .B(n459), .Y(n916) );
  XOR2X1 U764 ( .A(n616), .B(n609), .Y(n542) );
  XNOR2X1 U765 ( .A(n417), .B(n418), .Y(n416) );
  XOR2X1 U766 ( .A(n396), .B(n475), .Y(n321) );
  XOR2X1 U767 ( .A(n825), .B(n545), .Y(n614) );
  XOR2X1 U768 ( .A(n523), .B(n676), .Y(n288) );
  XOR2X1 U769 ( .A(n300), .B(n463), .Y(n683) );
  XOR2X1 U770 ( .A(n657), .B(n249), .Y(n654) );
  XOR2X1 U771 ( .A(n658), .B(n280), .Y(n657) );
  XOR2X1 U772 ( .A(n1410), .B(n249), .Y(n1403) );
  XOR2X1 U773 ( .A(n1028), .B(n270), .Y(n1410) );
  XOR2X1 U774 ( .A(n832), .B(n833), .Y(n456) );
  XOR2X1 U775 ( .A(n727), .B(n328), .Y(n724) );
  XOR2X1 U776 ( .A(n728), .B(n360), .Y(n727) );
  XOR2X1 U777 ( .A(n1175), .B(n328), .Y(n1169) );
  XOR2X1 U778 ( .A(n1163), .B(n350), .Y(n1175) );
  XOR2X1 U779 ( .A(n1126), .B(n756), .Y(n378) );
  XOR2X1 U780 ( .A(n372), .B(n1418), .Y(n1043) );
  XOR2X1 U781 ( .A(n584), .B(n489), .Y(n581) );
  XNOR2X1 U782 ( .A(n510), .B(n520), .Y(n584) );
  XOR2X1 U783 ( .A(n1255), .B(n409), .Y(n1249) );
  XOR2X1 U784 ( .A(n970), .B(n429), .Y(n1255) );
  XOR2X1 U785 ( .A(n801), .B(n409), .Y(n798) );
  XOR2X1 U786 ( .A(n802), .B(n439), .Y(n801) );
  XOR2X1 U787 ( .A(n1331), .B(n489), .Y(n1327) );
  XNOR2X1 U788 ( .A(n594), .B(n509), .Y(n1331) );
  XOR2X1 U789 ( .A(n697), .B(n1695), .Y(n1384) );
  XOR2X1 U790 ( .A(n1005), .B(n1006), .Y(n1003) );
  XOR2X1 U791 ( .A(n488), .B(n633), .Y(n1006) );
  XOR2X1 U792 ( .A(n1125), .B(n764), .Y(n1133) );
  XOR2X1 U793 ( .A(n763), .B(n764), .Y(n760) );
  XOR2X1 U794 ( .A(n765), .B(n393), .Y(n763) );
  XOR2X1 U795 ( .A(n1308), .B(n472), .Y(n1306) );
  XNOR2X1 U796 ( .A(n935), .B(n857), .Y(n1308) );
  XOR2X1 U797 ( .A(n843), .B(n844), .Y(n840) );
  XOR2X1 U798 ( .A(n845), .B(n1684), .Y(n843) );
  XOR2X1 U799 ( .A(n710), .B(n711), .Y(n707) );
  XOR2X1 U800 ( .A(n712), .B(n327), .Y(n711) );
  XOR2X1 U801 ( .A(n1302), .B(n926), .Y(n1295) );
  XNOR2X1 U802 ( .A(n834), .B(n472), .Y(n1302) );
  XOR2X1 U803 ( .A(n1377), .B(n557), .Y(n1371) );
  XNOR2X1 U804 ( .A(n546), .B(n999), .Y(n1377) );
  XNOR2X1 U805 ( .A(n310), .B(n1056), .Y(n1052) );
  XOR2X1 U806 ( .A(n535), .B(n463), .Y(n1056) );
  XOR2X1 U807 ( .A(n755), .B(n390), .Y(n1218) );
  XOR2X1 U808 ( .A(n1427), .B(n1064), .Y(n1453) );
  XNOR2X1 U809 ( .A(n392), .B(n756), .Y(n752) );
  XOR2X1 U810 ( .A(n981), .B(n982), .Y(n974) );
  XNOR2X1 U811 ( .A(n605), .B(n597), .Y(n981) );
  XOR2X1 U812 ( .A(n1357), .B(n532), .Y(n1349) );
  XOR2X1 U813 ( .A(n978), .B(n982), .Y(n1357) );
  XOR2X1 U814 ( .A(n327), .B(n774), .Y(n1142) );
  XNOR2X1 U815 ( .A(n1125), .B(n1126), .Y(n1207) );
  XOR2X1 U816 ( .A(n856), .B(n857), .Y(n849) );
  XOR2X1 U817 ( .A(n858), .B(n859), .Y(n856) );
  XOR2X1 U818 ( .A(n1202), .B(n1119), .Y(n1193) );
  XNOR2X1 U819 ( .A(n1114), .B(n1113), .Y(n1202) );
  XOR2X1 U820 ( .A(n567), .B(n568), .Y(n564) );
  XOR2X1 U821 ( .A(n569), .B(n488), .Y(n568) );
  XOR2X1 U822 ( .A(n310), .B(n311), .Y(n306) );
  XOR2X1 U823 ( .A(n497), .B(n575), .Y(n574) );
  XOR2X1 U824 ( .A(n518), .B(n519), .Y(n514) );
  XOR2X1 U825 ( .A(n520), .B(n1670), .Y(n518) );
  XOR2X1 U826 ( .A(n908), .B(n909), .Y(n902) );
  XNOR2X1 U827 ( .A(n910), .B(n822), .Y(n908) );
  XOR2X1 U828 ( .A(n1281), .B(n909), .Y(n1273) );
  XOR2X1 U829 ( .A(n1048), .B(n821), .Y(n1281) );
  XOR2X1 U830 ( .A(n896), .B(n897), .Y(n892) );
  XOR2X1 U831 ( .A(n429), .B(n1679), .Y(n896) );
  XOR2X1 U832 ( .A(n278), .B(n279), .Y(n274) );
  XOR2X1 U833 ( .A(n280), .B(n1657), .Y(n278) );
  XOR2X1 U834 ( .A(n746), .B(n371), .Y(n741) );
  XNOR2X1 U835 ( .A(n747), .B(n748), .Y(n746) );
  XNOR2X1 U836 ( .A(n519), .B(n592), .Y(n588) );
  XOR2X1 U837 ( .A(n593), .B(n594), .Y(n592) );
  XOR2X1 U838 ( .A(n1105), .B(n1106), .Y(n1101) );
  XOR2X1 U839 ( .A(n350), .B(n1691), .Y(n1105) );
  XNOR2X1 U840 ( .A(n968), .B(n1345), .Y(n1335) );
  XOR2X1 U841 ( .A(n593), .B(n510), .Y(n1345) );
  XNOR2X1 U842 ( .A(n834), .B(n835), .Y(n827) );
  XOR2X1 U843 ( .A(n836), .B(n471), .Y(n835) );
  XNOR2X1 U844 ( .A(n543), .B(n544), .Y(n537) );
  XOR2X1 U845 ( .A(n545), .B(n546), .Y(n544) );
  XNOR2X1 U846 ( .A(n624), .B(n998), .Y(n994) );
  XOR2X1 U847 ( .A(n543), .B(n999), .Y(n998) );
  XOR2X1 U848 ( .A(n437), .B(n438), .Y(n433) );
  XOR2X1 U849 ( .A(n439), .B(n1679), .Y(n437) );
  XOR2X1 U850 ( .A(n967), .B(n968), .Y(n963) );
  XOR2X1 U851 ( .A(n509), .B(n1670), .Y(n967) );
  XOR2X1 U852 ( .A(n358), .B(n359), .Y(n354) );
  XOR2X1 U853 ( .A(n360), .B(n1691), .Y(n358) );
  XOR2X1 U854 ( .A(n1656), .B(n1392), .Y(n1390) );
  XOR2X1 U855 ( .A(n251), .B(n404), .Y(n1392) );
  XOR2X1 U856 ( .A(n775), .B(n776), .Y(n770) );
  XOR2X1 U857 ( .A(n1689), .B(n777), .Y(n776) );
  XOR2X1 U858 ( .A(n702), .B(n1468), .Y(n1465) );
  XOR2X1 U859 ( .A(n243), .B(n484), .Y(n1468) );
  XNOR2X1 U860 ( .A(n300), .B(n301), .Y(n296) );
  XOR2X1 U861 ( .A(n302), .B(n1701), .Y(n301) );
  XOR2X1 U862 ( .A(n421), .B(n878), .Y(n875) );
  XOR2X1 U863 ( .A(n879), .B(n427), .Y(n878) );
  XOR2X1 U864 ( .A(n469), .B(n470), .Y(n465) );
  XOR2X1 U865 ( .A(n471), .B(n472), .Y(n470) );
  XOR2X1 U866 ( .A(n554), .B(n555), .Y(n550) );
  XOR2X1 U867 ( .A(n556), .B(n557), .Y(n555) );
  XOR2X1 U868 ( .A(n1671), .B(n959), .Y(n954) );
  XOR2X1 U869 ( .A(n520), .B(n594), .Y(n959) );
  XOR2X1 U870 ( .A(n927), .B(n1291), .Y(n1285) );
  XOR2X1 U871 ( .A(n832), .B(n845), .Y(n1291) );
  XOR2X1 U872 ( .A(n507), .B(n508), .Y(n505) );
  XOR2X1 U873 ( .A(n509), .B(n510), .Y(n508) );
  XOR2X1 U874 ( .A(n396), .B(n1073), .Y(n1069) );
  XOR2X1 U875 ( .A(n248), .B(n314), .Y(n1073) );
  XOR2X1 U876 ( .A(n262), .B(n1018), .Y(n1016) );
  XOR2X1 U877 ( .A(n251), .B(n268), .Y(n1018) );
  XOR2X1 U878 ( .A(n342), .B(n1087), .Y(n1084) );
  XOR2X1 U879 ( .A(n1088), .B(n348), .Y(n1087) );
  XOR2X1 U880 ( .A(n989), .B(n990), .Y(n986) );
  XOR2X1 U881 ( .A(n609), .B(n556), .Y(n990) );
  XOR2X1 U882 ( .A(n710), .B(n1230), .Y(n1227) );
  XOR2X1 U883 ( .A(n1694), .B(n775), .Y(n1230) );
  XOR2X1 U884 ( .A(n390), .B(n391), .Y(n386) );
  XOR2X1 U885 ( .A(n392), .B(n393), .Y(n391) );
  XOR2X1 U886 ( .A(n258), .B(n1660), .Y(n257) );
  XOR2X1 U887 ( .A(n641), .B(n1656), .Y(n640) );
  XOR2X1 U888 ( .A(n852), .B(n934), .Y(n931) );
  XOR2X1 U889 ( .A(n408), .B(n854), .Y(n934) );
  XOR2X1 U890 ( .A(n268), .B(n269), .Y(n266) );
  XOR2X1 U891 ( .A(n270), .B(n1658), .Y(n269) );
  XOR2X1 U892 ( .A(n1682), .B(n888), .Y(n883) );
  XOR2X1 U893 ( .A(n439), .B(n1678), .Y(n888) );
  XOR2X1 U894 ( .A(n427), .B(n428), .Y(n425) );
  XOR2X1 U895 ( .A(n429), .B(n1686), .Y(n428) );
  XOR2X1 U896 ( .A(n261), .B(n1027), .Y(n1022) );
  XOR2X1 U897 ( .A(n280), .B(n1664), .Y(n1027) );
  XOR2X1 U898 ( .A(n348), .B(n349), .Y(n346) );
  XOR2X1 U899 ( .A(n350), .B(n1692), .Y(n349) );
  XOR2X1 U900 ( .A(n341), .B(n1097), .Y(n1092) );
  XOR2X1 U901 ( .A(n360), .B(n1700), .Y(n1097) );
  XOR2X1 U902 ( .A(n1036), .B(n1661), .Y(n1032) );
  XOR2X1 U903 ( .A(n270), .B(n1657), .Y(n1036) );
  INVX1 U904 ( .A(n1163), .Y(n1700) );
  INVX1 U905 ( .A(n970), .Y(n1678) );
  INVX1 U906 ( .A(n1028), .Y(n1664) );
  INVX1 U907 ( .A(n1427), .Y(n1701) );
  INVX1 U908 ( .A(n765), .Y(n1688) );
  INVX1 U909 ( .A(n989), .Y(n1665) );
  INVX1 U910 ( .A(n927), .Y(n1680) );
  INVX1 U911 ( .A(n1048), .Y(n1683) );
  INVX1 U912 ( .A(n372), .Y(n1659) );
  INVX1 U913 ( .A(n978), .Y(n1672) );
  NOR2BX1 U914 ( .AN(n1477), .B(n1476), .Y(n242) );
  NAND2X1 U915 ( .A(n1478), .B(n1483), .Y(n1485) );
  NAND2X1 U916 ( .A(n1489), .B(n1469), .Y(n1483) );
  INVX1 U917 ( .A(n1489), .Y(n1706) );
  OA22X1 U918 ( .A0(n1631), .A1(n137), .B0(n1630), .B1(n90), .Y(n233) );
  OA22X1 U919 ( .A0(n1633), .A1(n146), .B0(n1629), .B1(n102), .Y(n210) );
  OA22X1 U920 ( .A0(n1632), .A1(n125), .B0(n1628), .B1(n79), .Y(n224) );
  OA22X1 U921 ( .A0(n1633), .A1(n114), .B0(n1629), .B1(n65), .Y(n216) );
  OA22X1 U922 ( .A0(n1632), .A1(n126), .B0(n1628), .B1(n80), .Y(n226) );
  OA22X1 U923 ( .A0(n1633), .A1(n117), .B0(n1629), .B1(n67), .Y(n217) );
  OA22X1 U924 ( .A0(n1633), .A1(n148), .B0(n1629), .B1(n103), .Y(n211) );
  OA22X1 U925 ( .A0(n1631), .A1(n138), .B0(n205), .B1(n92), .Y(n234) );
  NOR2X1 U926 ( .A(n1709), .B(n1710), .Y(n1475) );
  NOR2X1 U927 ( .A(n1), .B(n8), .Y(n1709) );
  NOR2X1 U928 ( .A(n1705), .B(n1707), .Y(n1710) );
  NOR2X1 U929 ( .A(n8), .B(n7), .Y(n1477) );
  NAND3X1 U930 ( .A(n57), .B(n56), .C(n860), .Y(n202) );
  OR4X1 U931 ( .A(round[0]), .B(round[1]), .C(round[2]), .D(round[3]), .Y(
        n1476) );
  OAI221XL U932 ( .A0(n1639), .A1(n32), .B0(n1635), .B1(n176), .C0(n227), .Y(
        tmp_sboxw[18]) );
  OA22X1 U933 ( .A0(n1632), .A1(n127), .B0(n1628), .B1(n81), .Y(n227) );
  OAI221XL U934 ( .A0(n1638), .A1(n51), .B0(n1636), .B1(n197), .C0(n214), .Y(
        tmp_sboxw[2]) );
  OA22X1 U935 ( .A0(n1633), .A1(n149), .B0(n1629), .B1(n104), .Y(n214) );
  OAI221XL U936 ( .A0(n1639), .A1(n22), .B0(n1635), .B1(n161), .C0(n218), .Y(
        tmp_sboxw[26]) );
  OA22X1 U937 ( .A0(n1632), .A1(n118), .B0(n1628), .B1(n68), .Y(n218) );
  OAI221XL U938 ( .A0(n1637), .A1(n43), .B0(n1634), .B1(n185), .C0(n235), .Y(
        tmp_sboxw[10]) );
  OA22X1 U939 ( .A0(n1631), .A1(n139), .B0(n205), .B1(n93), .Y(n235) );
  OA22X1 U940 ( .A0(n1631), .A1(n130), .B0(n205), .B1(n84), .Y(n229) );
  OA22X1 U941 ( .A0(n1631), .A1(n151), .B0(n205), .B1(n106), .Y(n236) );
  OA22X1 U942 ( .A0(n204), .A1(n140), .B0(n1630), .B1(n94), .Y(n203) );
  OA22X1 U943 ( .A0(n1632), .A1(n119), .B0(n1628), .B1(n69), .Y(n219) );
  OA22X1 U944 ( .A0(n1632), .A1(n121), .B0(n1628), .B1(n70), .Y(n220) );
  OA22X1 U945 ( .A0(n1631), .A1(n129), .B0(n205), .B1(n83), .Y(n228) );
  OA22X1 U946 ( .A0(n204), .A1(n141), .B0(n1630), .B1(n95), .Y(n206) );
  OA22X1 U947 ( .A0(n1632), .A1(n150), .B0(n1628), .B1(n105), .Y(n225) );
  OAI221XL U948 ( .A0(n292), .A1(n192), .B0(n161), .B1(n2), .C0(n293), .Y(
        n1496) );
  XNOR2X1 U949 ( .A(round_key[122]), .B(block[122]), .Y(n292) );
  AOI222XL U950 ( .A0(new_sboxw[26]), .A1(n156), .B0(n108), .B1(n294), .C0(n82), .C1(n295), .Y(n293) );
  XOR2X1 U951 ( .A(n296), .B(n297), .Y(n295) );
  OAI221XL U952 ( .A0(n547), .A1(n239), .B0(n198), .B1(n160), .C0(n548), .Y(
        n1521) );
  XNOR2X1 U953 ( .A(round_key[65]), .B(block[65]), .Y(n547) );
  AOI222XL U954 ( .A0(new_sboxw[1]), .A1(n153), .B0(n131), .B1(n310), .C0(n91), 
        .C1(n549), .Y(n548) );
  XOR2X1 U955 ( .A(n550), .B(n551), .Y(n549) );
  OAI221XL U956 ( .A0(n617), .A1(n239), .B0(n119), .B1(n60), .C0(n618), .Y(
        n1528) );
  XNOR2X1 U957 ( .A(round_key[89]), .B(block[89]), .Y(n617) );
  AOI222XL U958 ( .A0(n33), .A1(new_sboxw[25]), .B0(n101), .B1(n543), .C0(n96), 
        .C1(n619), .Y(n618) );
  XOR2X1 U959 ( .A(n620), .B(n621), .Y(n619) );
  OAI221XL U960 ( .A0(n686), .A1(n190), .B0(n129), .B1(n59), .C0(n687), .Y(
        n1536) );
  XNOR2X1 U961 ( .A(round_key[113]), .B(block[113]), .Y(n686) );
  AOI222XL U962 ( .A0(n36), .A1(new_sboxw[17]), .B0(n131), .B1(n1665), .C0(n78), .C1(n688), .Y(n687) );
  XOR2X1 U963 ( .A(n689), .B(n690), .Y(n688) );
  OAI221XL U964 ( .A0(n626), .A1(n743), .B0(n121), .B1(n60), .C0(n627), .Y(
        n1529) );
  XNOR2X1 U965 ( .A(round_key[88]), .B(block[88]), .Y(n626) );
  AOI222XL U966 ( .A0(n33), .A1(new_sboxw[24]), .B0(n135), .B1(n1695), .C0(n88), .C1(n628), .Y(n627) );
  XOR2X1 U967 ( .A(n629), .B(n630), .Y(n628) );
  OAI221XL U968 ( .A0(n695), .A1(n190), .B0(n130), .B1(n59), .C0(n696), .Y(
        n1537) );
  XNOR2X1 U969 ( .A(round_key[112]), .B(block[112]), .Y(n695) );
  AOI222XL U970 ( .A0(n36), .A1(new_sboxw[16]), .B0(n101), .B1(n697), .C0(n78), 
        .C1(n698), .Y(n696) );
  XOR2X1 U971 ( .A(n699), .B(n700), .Y(n698) );
  OAI221XL U972 ( .A0(n473), .A1(n194), .B0(n187), .B1(n160), .C0(n474), .Y(
        n1514) );
  XNOR2X1 U973 ( .A(round_key[40]), .B(block[40]), .Y(n473) );
  AOI222XL U974 ( .A0(new_sboxw[8]), .A1(n153), .B0(n101), .B1(n475), .C0(n85), 
        .C1(n476), .Y(n474) );
  XOR2X1 U975 ( .A(n477), .B(n478), .Y(n476) );
  OAI221XL U976 ( .A0(n928), .A1(n174), .B0(n70), .B1(n25), .C0(n929), .Y(
        n1561) );
  XNOR2X1 U977 ( .A(round_key[56]), .B(block[56]), .Y(n928) );
  AOI222XL U978 ( .A0(n17), .A1(new_sboxw[24]), .B0(n107), .B1(n853), .C0(n74), 
        .C1(n930), .Y(n929) );
  XOR2X1 U979 ( .A(n931), .B(n932), .Y(n930) );
  OAI221XL U980 ( .A0(n704), .A1(n190), .B0(n132), .B1(n59), .C0(n705), .Y(
        n1538) );
  XNOR2X1 U981 ( .A(round_key[15]), .B(block[15]), .Y(n704) );
  AOI222XL U982 ( .A0(n36), .A1(new_sboxw[15]), .B0(n131), .B1(n1666), .C0(n78), .C1(n706), .Y(n705) );
  XOR2X1 U983 ( .A(n707), .B(n708), .Y(n706) );
  OAI221XL U984 ( .A0(n951), .A1(n174), .B0(n76), .B1(n25), .C0(n952), .Y(
        n1564) );
  XNOR2X1 U985 ( .A(round_key[85]), .B(block[85]), .Y(n951) );
  AOI222XL U986 ( .A0(n17), .A1(new_sboxw[21]), .B0(n107), .B1(n1675), .C0(n74), .C1(n953), .Y(n952) );
  XOR2X1 U987 ( .A(n954), .B(n506), .Y(n953) );
  OAI221XL U988 ( .A0(n253), .A1(n192), .B0(n154), .B1(n165), .C0(n254), .Y(
        n1492) );
  XNOR2X1 U989 ( .A(round_key[126]), .B(block[126]), .Y(n253) );
  AOI222XL U990 ( .A0(new_sboxw[30]), .A1(n241), .B0(n108), .B1(n251), .C0(n82), .C1(n255), .Y(n254) );
  XOR2X1 U991 ( .A(n256), .B(n257), .Y(n255) );
  OAI221XL U992 ( .A0(n263), .A1(n192), .B0(n157), .B1(n165), .C0(n264), .Y(
        n1493) );
  XNOR2X1 U993 ( .A(round_key[125]), .B(block[125]), .Y(n263) );
  AOI222XL U994 ( .A0(new_sboxw[29]), .A1(n156), .B0(n108), .B1(n261), .C0(n82), .C1(n265), .Y(n264) );
  XOR2X1 U995 ( .A(n266), .B(n267), .Y(n265) );
  OAI221XL U996 ( .A0(n1007), .A1(n172), .B0(n86), .B1(n19), .C0(n1008), .Y(
        n1570) );
  XNOR2X1 U997 ( .A(round_key[111]), .B(block[111]), .Y(n1007) );
  AOI222XL U998 ( .A0(n15), .A1(new_sboxw[15]), .B0(n242), .B1(n1681), .C0(n72), .C1(n1009), .Y(n1008) );
  XOR2X1 U999 ( .A(n1010), .B(n1011), .Y(n1009) );
  OAI221XL U1000 ( .A0(n570), .A1(n192), .B0(n110), .B1(n559), .C0(n571), .Y(
        n1523) );
  XNOR2X1 U1001 ( .A(round_key[94]), .B(block[94]), .Y(n570) );
  AOI222XL U1002 ( .A0(n36), .A1(new_sboxw[30]), .B0(n131), .B1(n569), .C0(n88), .C1(n572), .Y(n571) );
  XOR2X1 U1003 ( .A(n573), .B(n574), .Y(n572) );
  OAI221XL U1004 ( .A0(n502), .A1(n194), .B0(n193), .B1(n160), .C0(n503), .Y(
        n1517) );
  XNOR2X1 U1005 ( .A(round_key[69]), .B(block[69]), .Y(n502) );
  AOI222XL U1006 ( .A0(new_sboxw[5]), .A1(n153), .B0(n133), .B1(n1663), .C0(
        n91), .C1(n504), .Y(n503) );
  XOR2X1 U1007 ( .A(n505), .B(n506), .Y(n504) );
  OAI221XL U1008 ( .A0(n651), .A1(n190), .B0(n124), .B1(n60), .C0(n652), .Y(
        n1532) );
  XNOR2X1 U1009 ( .A(round_key[117]), .B(block[117]), .Y(n651) );
  AOI222XL U1010 ( .A0(n33), .A1(new_sboxw[21]), .B0(n135), .B1(n507), .C0(n78), .C1(n653), .Y(n652) );
  XOR2X1 U1011 ( .A(n654), .B(n655), .Y(n653) );
  OAI221XL U1012 ( .A0(n430), .A1(n239), .B0(n183), .B1(n162), .C0(n431), .Y(
        n1510) );
  XNOR2X1 U1013 ( .A(round_key[44]), .B(block[44]), .Y(n430) );
  AOI222XL U1014 ( .A0(new_sboxw[12]), .A1(n155), .B0(n133), .B1(n280), .C0(
        n85), .C1(n432), .Y(n431) );
  XOR2X1 U1015 ( .A(n433), .B(n434), .Y(n432) );
  OAI221XL U1016 ( .A0(n880), .A1(n180), .B0(n63), .B1(n864), .C0(n881), .Y(
        n1556) );
  XNOR2X1 U1017 ( .A(round_key[61]), .B(block[61]), .Y(n880) );
  AOI222XL U1018 ( .A0(n17), .A1(new_sboxw[29]), .B0(n115), .B1(n427), .C0(n75), .C1(n882), .Y(n881) );
  XOR2X1 U1019 ( .A(n883), .B(n426), .Y(n882) );
  OAI221XL U1020 ( .A0(n644), .A1(n190), .B0(n123), .B1(n60), .C0(n645), .Y(
        n1531) );
  XNOR2X1 U1021 ( .A(round_key[118]), .B(block[118]), .Y(n644) );
  AOI222XL U1022 ( .A0(n33), .A1(new_sboxw[22]), .B0(n144), .B1(n498), .C0(n78), .C1(n646), .Y(n645) );
  XOR2X1 U1023 ( .A(n647), .B(n648), .Y(n646) );
  OAI221XL U1024 ( .A0(n595), .A1(n743), .B0(n117), .B1(n60), .C0(n596), .Y(
        n1526) );
  XNOR2X1 U1025 ( .A(round_key[91]), .B(block[91]), .Y(n595) );
  AOI222XL U1026 ( .A0(n33), .A1(new_sboxw[27]), .B0(n101), .B1(n597), .C0(n88), .C1(n598), .Y(n596) );
  XOR2X1 U1027 ( .A(n599), .B(n600), .Y(n598) );
  OAI221XL U1028 ( .A0(n677), .A1(n190), .B0(n127), .B1(n59), .C0(n678), .Y(
        n1535) );
  XNOR2X1 U1029 ( .A(round_key[114]), .B(block[114]), .Y(n677) );
  AOI222XL U1030 ( .A0(n36), .A1(new_sboxw[18]), .B0(n101), .B1(n616), .C0(n78), .C1(n679), .Y(n678) );
  XOR2X1 U1031 ( .A(n680), .B(n681), .Y(n679) );
  OAI221XL U1032 ( .A0(n450), .A1(n239), .B0(n185), .B1(n162), .C0(n451), .Y(
        n1512) );
  XNOR2X1 U1033 ( .A(round_key[42]), .B(block[42]), .Y(n450) );
  AOI222XL U1034 ( .A0(new_sboxw[10]), .A1(n155), .B0(n144), .B1(n452), .C0(
        n88), .C1(n453), .Y(n451) );
  XOR2X1 U1035 ( .A(n454), .B(n455), .Y(n453) );
  OAI221XL U1036 ( .A0(n1066), .A1(n172), .B0(n95), .B1(n18), .C0(n1067), .Y(
        n1577) );
  XNOR2X1 U1037 ( .A(round_key[104]), .B(block[104]), .Y(n1066) );
  AOI222XL U1038 ( .A0(n14), .A1(new_sboxw[8]), .B0(n242), .B1(n854), .C0(n72), 
        .C1(n1068), .Y(n1067) );
  XOR2X1 U1039 ( .A(n1069), .B(n1070), .Y(n1068) );
  OAI221XL U1040 ( .A0(n422), .A1(n194), .B0(n182), .B1(n162), .C0(n423), .Y(
        n1509) );
  XNOR2X1 U1041 ( .A(round_key[45]), .B(block[45]), .Y(n422) );
  AOI222XL U1042 ( .A0(new_sboxw[13]), .A1(n155), .B0(n131), .B1(n268), .C0(
        n96), .C1(n424), .Y(n423) );
  XOR2X1 U1043 ( .A(n425), .B(n426), .Y(n424) );
  OAI221XL U1044 ( .A0(n1029), .A1(n172), .B0(n90), .B1(n19), .C0(n1030), .Y(
        n1573) );
  XNOR2X1 U1045 ( .A(round_key[108]), .B(block[108]), .Y(n1029) );
  AOI222XL U1046 ( .A0(n15), .A1(new_sboxw[12]), .B0(n107), .B1(n429), .C0(n72), .C1(n1031), .Y(n1030) );
  XOR2X1 U1047 ( .A(n1032), .B(n1033), .Y(n1031) );
  OAI221XL U1048 ( .A0(n461), .A1(n743), .B0(n186), .B1(n162), .C0(n462), .Y(
        n1513) );
  XNOR2X1 U1049 ( .A(round_key[41]), .B(block[41]), .Y(n461) );
  AOI222XL U1050 ( .A0(new_sboxw[9]), .A1(n153), .B0(n135), .B1(n463), .C0(n85), .C1(n464), .Y(n462) );
  XOR2X1 U1051 ( .A(n465), .B(n466), .Y(n464) );
  OAI221XL U1052 ( .A0(n991), .A1(n174), .B0(n83), .B1(n19), .C0(n992), .Y(
        n1568) );
  XNOR2X1 U1053 ( .A(round_key[81]), .B(block[81]), .Y(n991) );
  AOI222XL U1054 ( .A0(n15), .A1(new_sboxw[17]), .B0(n242), .B1(n1680), .C0(
        n74), .C1(n993), .Y(n992) );
  XOR2X1 U1055 ( .A(n994), .B(n995), .Y(n993) );
  OAI221XL U1056 ( .A0(n786), .A1(n189), .B0(n143), .B1(n40), .C0(n787), .Y(
        n1547) );
  XNOR2X1 U1057 ( .A(round_key[38]), .B(block[38]), .Y(n786) );
  AOI222XL U1058 ( .A0(n30), .A1(new_sboxw[6]), .B0(n113), .B1(n788), .C0(n77), 
        .C1(n789), .Y(n787) );
  XOR2X1 U1059 ( .A(n790), .B(n791), .Y(n789) );
  OAI221XL U1060 ( .A0(n812), .A1(n180), .B0(n148), .B1(n40), .C0(n813), .Y(
        n1550) );
  XNOR2X1 U1061 ( .A(round_key[35]), .B(block[35]), .Y(n812) );
  AOI222XL U1062 ( .A0(n30), .A1(new_sboxw[3]), .B0(n115), .B1(n1672), .C0(n75), .C1(n814), .Y(n813) );
  XOR2X1 U1063 ( .A(n815), .B(n816), .Y(n814) );
  OAI221XL U1064 ( .A0(n1393), .A1(n1486), .B0(n47), .B1(n9), .C0(n1394), .Y(
        n1611) );
  XNOR2X1 U1065 ( .A(round_key[102]), .B(block[102]), .Y(n1393) );
  AOI222XL U1066 ( .A0(n4), .A1(new_sboxw[6]), .B0(n128), .B1(n338), .C0(n97), 
        .C1(n1395), .Y(n1394) );
  XOR2X1 U1067 ( .A(n1396), .B(n1397), .Y(n1395) );
  OAI221XL U1068 ( .A0(n281), .A1(n192), .B0(n159), .B1(n2), .C0(n282), .Y(
        n1495) );
  XNOR2X1 U1069 ( .A(round_key[123]), .B(block[123]), .Y(n281) );
  AOI222XL U1070 ( .A0(new_sboxw[27]), .A1(n156), .B0(n108), .B1(n283), .C0(
        n82), .C1(n284), .Y(n282) );
  XOR2X1 U1071 ( .A(n285), .B(n286), .Y(n284) );
  OAI221XL U1072 ( .A0(n440), .A1(n200), .B0(n184), .B1(n162), .C0(n441), .Y(
        n1511) );
  XNOR2X1 U1073 ( .A(round_key[43]), .B(block[43]), .Y(n440) );
  AOI222XL U1074 ( .A0(new_sboxw[11]), .A1(n155), .B0(n133), .B1(n442), .C0(
        n96), .C1(n443), .Y(n441) );
  XOR2X1 U1075 ( .A(n444), .B(n445), .Y(n443) );
  OAI221XL U1076 ( .A0(n1013), .A1(n172), .B0(n87), .B1(n19), .C0(n1014), .Y(
        n1571) );
  XNOR2X1 U1077 ( .A(round_key[110]), .B(block[110]), .Y(n1013) );
  AOI222XL U1078 ( .A0(n15), .A1(new_sboxw[14]), .B0(n135), .B1(n879), .C0(n72), .C1(n1015), .Y(n1014) );
  XOR2X1 U1079 ( .A(n1016), .B(n1017), .Y(n1015) );
  OAI221XL U1080 ( .A0(n331), .A1(n239), .B0(n168), .B1(n165), .C0(n332), .Y(
        n1500) );
  XNOR2X1 U1081 ( .A(round_key[22]), .B(block[22]), .Y(n331) );
  AOI222XL U1082 ( .A0(new_sboxw[22]), .A1(n156), .B0(n111), .B1(n333), .C0(
        n91), .C1(n334), .Y(n332) );
  XOR2X1 U1083 ( .A(n335), .B(n336), .Y(n334) );
  OAI221XL U1084 ( .A0(n1315), .A1(n166), .B0(n38), .B1(n10), .C0(n1316), .Y(
        n1603) );
  XNOR2X1 U1085 ( .A(round_key[78]), .B(block[78]), .Y(n1315) );
  AOI222XL U1086 ( .A0(n5), .A1(new_sboxw[14]), .B0(n120), .B1(n712), .C0(n61), 
        .C1(n1317), .Y(n1316) );
  XOR2X1 U1087 ( .A(n1318), .B(n1319), .Y(n1317) );
  OAI221XL U1088 ( .A0(n837), .A1(n180), .B0(n150), .B1(n40), .C0(n838), .Y(
        n1552) );
  XNOR2X1 U1089 ( .A(round_key[33]), .B(block[33]), .Y(n837) );
  AOI222XL U1090 ( .A0(n30), .A1(new_sboxw[1]), .B0(n115), .B1(n546), .C0(n75), 
        .C1(n839), .Y(n838) );
  XOR2X1 U1091 ( .A(n840), .B(n841), .Y(n839) );
  OAI221XL U1092 ( .A0(n412), .A1(n743), .B0(n181), .B1(n162), .C0(n413), .Y(
        n1508) );
  XNOR2X1 U1093 ( .A(round_key[46]), .B(block[46]), .Y(n412) );
  AOI222XL U1094 ( .A0(new_sboxw[14]), .A1(n155), .B0(n111), .B1(n1660), .C0(
        n88), .C1(n414), .Y(n413) );
  XOR2X1 U1095 ( .A(n415), .B(n416), .Y(n414) );
  OAI221XL U1096 ( .A0(n872), .A1(n180), .B0(n62), .B1(n864), .C0(n873), .Y(
        n1555) );
  XNOR2X1 U1097 ( .A(round_key[62]), .B(block[62]), .Y(n872) );
  AOI222XL U1098 ( .A0(n866), .A1(new_sboxw[30]), .B0(n115), .B1(n417), .C0(
        n75), .C1(n874), .Y(n873) );
  XOR2X1 U1099 ( .A(n875), .B(n876), .Y(n874) );
  OAI221XL U1100 ( .A0(n1081), .A1(n172), .B0(n99), .B1(n18), .C0(n1082), .Y(
        n1579) );
  XNOR2X1 U1101 ( .A(round_key[6]), .B(block[6]), .Y(n1081) );
  AOI222XL U1102 ( .A0(n14), .A1(new_sboxw[6]), .B0(n133), .B1(n785), .C0(n72), 
        .C1(n1083), .Y(n1082) );
  XOR2X1 U1103 ( .A(n1084), .B(n1085), .Y(n1083) );
  OAI221XL U1104 ( .A0(n521), .A1(n194), .B0(n196), .B1(n160), .C0(n522), .Y(
        n1519) );
  XNOR2X1 U1105 ( .A(round_key[67]), .B(block[67]), .Y(n521) );
  AOI222XL U1106 ( .A0(new_sboxw[3]), .A1(n153), .B0(n133), .B1(n523), .C0(n96), .C1(n524), .Y(n522) );
  XOR2X1 U1107 ( .A(n525), .B(n526), .Y(n524) );
  OAI221XL U1108 ( .A0(n668), .A1(n190), .B0(n126), .B1(n60), .C0(n669), .Y(
        n1534) );
  XNOR2X1 U1109 ( .A(round_key[115]), .B(block[115]), .Y(n668) );
  AOI222XL U1110 ( .A0(n36), .A1(new_sboxw[19]), .B0(n133), .B1(n604), .C0(n78), .C1(n670), .Y(n669) );
  XOR2X1 U1111 ( .A(n671), .B(n672), .Y(n670) );
  OAI221XL U1112 ( .A0(n312), .A1(n192), .B0(n164), .B1(n165), .C0(n313), .Y(
        n1498) );
  XNOR2X1 U1113 ( .A(round_key[120]), .B(block[120]), .Y(n312) );
  AOI222XL U1114 ( .A0(new_sboxw[24]), .A1(n156), .B0(n108), .B1(n314), .C0(
        n82), .C1(n315), .Y(n313) );
  XOR2X1 U1115 ( .A(n316), .B(n317), .Y(n315) );
  OAI221XL U1116 ( .A0(n394), .A1(n743), .B0(n178), .B1(n162), .C0(n395), .Y(
        n1506) );
  XNOR2X1 U1117 ( .A(round_key[16]), .B(block[16]), .Y(n394) );
  AOI222XL U1118 ( .A0(new_sboxw[16]), .A1(n155), .B0(n111), .B1(n396), .C0(
        n91), .C1(n397), .Y(n395) );
  XNOR2X1 U1119 ( .A(n398), .B(n399), .Y(n397) );
  OAI221XL U1120 ( .A0(n1309), .A1(n166), .B0(n37), .B1(n10), .C0(n1310), .Y(
        n1602) );
  XNOR2X1 U1121 ( .A(round_key[79]), .B(block[79]), .Y(n1309) );
  AOI222XL U1122 ( .A0(n5), .A1(new_sboxw[15]), .B0(n120), .B1(n1689), .C0(n61), .C1(n1311), .Y(n1310) );
  XOR2X1 U1123 ( .A(n1312), .B(n1313), .Y(n1311) );
  OAI221XL U1124 ( .A0(n899), .A1(n180), .B0(n67), .B1(n25), .C0(n900), .Y(
        n1558) );
  XNOR2X1 U1125 ( .A(round_key[59]), .B(block[59]), .Y(n899) );
  AOI222XL U1126 ( .A0(n17), .A1(new_sboxw[27]), .B0(n107), .B1(n821), .C0(n75), .C1(n901), .Y(n900) );
  XOR2X1 U1127 ( .A(n902), .B(n903), .Y(n901) );
  OAI221XL U1128 ( .A0(n971), .A1(n174), .B0(n80), .B1(n25), .C0(n972), .Y(
        n1566) );
  XNOR2X1 U1129 ( .A(round_key[83]), .B(block[83]), .Y(n971) );
  AOI222XL U1130 ( .A0(n15), .A1(new_sboxw[19]), .B0(n107), .B1(n822), .C0(n74), .C1(n973), .Y(n972) );
  XOR2X1 U1131 ( .A(n974), .B(n975), .Y(n973) );
  OAI221XL U1132 ( .A0(n578), .A1(n239), .B0(n112), .B1(n559), .C0(n579), .Y(
        n1524) );
  XNOR2X1 U1133 ( .A(round_key[93]), .B(block[93]), .Y(n578) );
  AOI222XL U1134 ( .A0(n33), .A1(new_sboxw[29]), .B0(n133), .B1(n497), .C0(n88), .C1(n580), .Y(n579) );
  XOR2X1 U1135 ( .A(n581), .B(n582), .Y(n580) );
  OAI221XL U1136 ( .A0(n823), .A1(n180), .B0(n149), .B1(n40), .C0(n824), .Y(
        n1551) );
  XNOR2X1 U1137 ( .A(round_key[34]), .B(block[34]), .Y(n823) );
  AOI222XL U1138 ( .A0(n30), .A1(new_sboxw[2]), .B0(n115), .B1(n825), .C0(n75), 
        .C1(n826), .Y(n824) );
  XOR2X1 U1139 ( .A(n827), .B(n828), .Y(n826) );
  OAI221XL U1140 ( .A0(n1049), .A1(n172), .B0(n93), .B1(n19), .C0(n1050), .Y(
        n1575) );
  XNOR2X1 U1141 ( .A(round_key[106]), .B(block[106]), .Y(n1049) );
  AOI222XL U1142 ( .A0(n15), .A1(new_sboxw[10]), .B0(n242), .B1(n836), .C0(n72), .C1(n1051), .Y(n1050) );
  XOR2X1 U1143 ( .A(n1052), .B(n1053), .Y(n1051) );
  OAI221XL U1144 ( .A0(n373), .A1(n194), .B0(n176), .B1(n162), .C0(n374), .Y(
        n1504) );
  XNOR2X1 U1145 ( .A(round_key[18]), .B(block[18]), .Y(n373) );
  AOI222XL U1146 ( .A0(new_sboxw[18]), .A1(n155), .B0(n111), .B1(n302), .C0(
        n96), .C1(n375), .Y(n374) );
  XOR2X1 U1147 ( .A(n376), .B(n377), .Y(n375) );
  OAI221XL U1148 ( .A0(n402), .A1(n200), .B0(n179), .B1(n162), .C0(n403), .Y(
        n1507) );
  XNOR2X1 U1149 ( .A(round_key[47]), .B(block[47]), .Y(n402) );
  AOI222XL U1150 ( .A0(new_sboxw[15]), .A1(n155), .B0(n111), .B1(n404), .C0(
        n82), .C1(n405), .Y(n403) );
  XOR2X1 U1151 ( .A(n406), .B(n407), .Y(n405) );
  OAI221XL U1152 ( .A0(n918), .A1(n174), .B0(n69), .B1(n25), .C0(n919), .Y(
        n1560) );
  XNOR2X1 U1153 ( .A(round_key[57]), .B(block[57]), .Y(n918) );
  AOI222XL U1154 ( .A0(n17), .A1(new_sboxw[25]), .B0(n107), .B1(n834), .C0(n74), .C1(n920), .Y(n919) );
  XOR2X1 U1155 ( .A(n921), .B(n922), .Y(n920) );
  OAI221XL U1156 ( .A0(n1378), .A1(n166), .B0(n45), .B1(n9), .C0(n1379), .Y(
        n1609) );
  XNOR2X1 U1157 ( .A(round_key[72]), .B(block[72]), .Y(n1378) );
  AOI222XL U1158 ( .A0(n4), .A1(new_sboxw[8]), .B0(n128), .B1(n1147), .C0(n61), 
        .C1(n1380), .Y(n1379) );
  XOR2X1 U1159 ( .A(n1381), .B(n1382), .Y(n1380) );
  OAI221XL U1160 ( .A0(n846), .A1(n180), .B0(n151), .B1(n40), .C0(n847), .Y(
        n1553) );
  XNOR2X1 U1161 ( .A(round_key[32]), .B(block[32]), .Y(n846) );
  AOI222XL U1162 ( .A0(new_sboxw[0]), .A1(n30), .B0(n115), .B1(n633), .C0(n75), 
        .C1(n848), .Y(n847) );
  XOR2X1 U1163 ( .A(n849), .B(n850), .Y(n848) );
  OAI221XL U1164 ( .A0(n1019), .A1(n172), .B0(n89), .B1(n19), .C0(n1020), .Y(
        n1572) );
  XNOR2X1 U1165 ( .A(round_key[109]), .B(block[109]), .Y(n1019) );
  AOI222XL U1166 ( .A0(n15), .A1(new_sboxw[13]), .B0(n242), .B1(n1682), .C0(
        n72), .C1(n1021), .Y(n1020) );
  XOR2X1 U1167 ( .A(n1022), .B(n267), .Y(n1021) );
  OAI221XL U1168 ( .A0(n343), .A1(n194), .B0(n169), .B1(n165), .C0(n344), .Y(
        n1501) );
  XNOR2X1 U1169 ( .A(round_key[21]), .B(block[21]), .Y(n343) );
  AOI222XL U1170 ( .A0(new_sboxw[21]), .A1(n156), .B0(n111), .B1(n258), .C0(
        n88), .C1(n345), .Y(n344) );
  XOR2X1 U1171 ( .A(n346), .B(n347), .Y(n345) );
  OAI221XL U1172 ( .A0(n1238), .A1(n170), .B0(n27), .B1(n12), .C0(n1239), .Y(
        n1595) );
  XNOR2X1 U1173 ( .A(round_key[54]), .B(block[54]), .Y(n1238) );
  AOI222XL U1174 ( .A0(n6), .A1(new_sboxw[22]), .B0(n116), .B1(n1088), .C0(n64), .C1(n1240), .Y(n1239) );
  XOR2X1 U1175 ( .A(n1241), .B(n1242), .Y(n1240) );
  OAI221XL U1176 ( .A0(n1038), .A1(n172), .B0(n92), .B1(n19), .C0(n1039), .Y(
        n1574) );
  XNOR2X1 U1177 ( .A(round_key[107]), .B(block[107]), .Y(n1038) );
  AOI222XL U1178 ( .A0(n15), .A1(new_sboxw[11]), .B0(n242), .B1(n1683), .C0(
        n72), .C1(n1040), .Y(n1039) );
  XOR2X1 U1179 ( .A(n1041), .B(n1042), .Y(n1040) );
  OAI221XL U1180 ( .A0(n303), .A1(n192), .B0(n163), .B1(n2), .C0(n304), .Y(
        n1497) );
  XNOR2X1 U1181 ( .A(round_key[121]), .B(block[121]), .Y(n303) );
  AOI222XL U1182 ( .A0(new_sboxw[25]), .A1(n156), .B0(n108), .B1(n1701), .C0(
        n82), .C1(n305), .Y(n304) );
  XOR2X1 U1183 ( .A(n306), .B(n307), .Y(n305) );
  OAI221XL U1184 ( .A0(n383), .A1(n239), .B0(n177), .B1(n162), .C0(n384), .Y(
        n1505) );
  XNOR2X1 U1185 ( .A(round_key[17]), .B(block[17]), .Y(n383) );
  AOI222XL U1186 ( .A0(new_sboxw[17]), .A1(n155), .B0(n111), .B1(n300), .C0(
        n91), .C1(n385), .Y(n384) );
  XOR2X1 U1187 ( .A(n386), .B(n387), .Y(n385) );
  OAI221XL U1188 ( .A0(n1089), .A1(n171), .B0(n100), .B1(n18), .C0(n1090), .Y(
        n1580) );
  XNOR2X1 U1189 ( .A(round_key[5]), .B(block[5]), .Y(n1089) );
  AOI222XL U1190 ( .A0(n14), .A1(new_sboxw[5]), .B0(n144), .B1(n418), .C0(n66), 
        .C1(n1091), .Y(n1090) );
  XOR2X1 U1191 ( .A(n1092), .B(n347), .Y(n1091) );
  OAI221XL U1192 ( .A0(n533), .A1(n743), .B0(n197), .B1(n160), .C0(n534), .Y(
        n1520) );
  XNOR2X1 U1193 ( .A(round_key[66]), .B(block[66]), .Y(n533) );
  AOI222XL U1194 ( .A0(new_sboxw[2]), .A1(n153), .B0(n101), .B1(n535), .C0(n91), .C1(n536), .Y(n534) );
  XOR2X1 U1195 ( .A(n537), .B(n538), .Y(n536) );
  OAI221XL U1196 ( .A0(n607), .A1(n200), .B0(n118), .B1(n60), .C0(n608), .Y(
        n1527) );
  XNOR2X1 U1197 ( .A(round_key[90]), .B(block[90]), .Y(n607) );
  AOI222XL U1198 ( .A0(n33), .A1(new_sboxw[26]), .B0(n133), .B1(n609), .C0(n96), .C1(n610), .Y(n608) );
  XOR2X1 U1199 ( .A(n611), .B(n612), .Y(n610) );
  OAI221XL U1200 ( .A0(n766), .A1(n189), .B0(n141), .B1(n40), .C0(n767), .Y(
        n1545) );
  XNOR2X1 U1201 ( .A(round_key[8]), .B(block[8]), .Y(n766) );
  AOI222XL U1202 ( .A0(n30), .A1(new_sboxw[8]), .B0(n113), .B1(n768), .C0(n77), 
        .C1(n769), .Y(n767) );
  XOR2X1 U1203 ( .A(n770), .B(n771), .Y(n769) );
  OAI221XL U1204 ( .A0(n911), .A1(n180), .B0(n68), .B1(n25), .C0(n912), .Y(
        n1559) );
  XNOR2X1 U1205 ( .A(round_key[58]), .B(block[58]), .Y(n911) );
  AOI222XL U1206 ( .A0(n17), .A1(new_sboxw[26]), .B0(n107), .B1(n832), .C0(n75), .C1(n913), .Y(n912) );
  XOR2X1 U1207 ( .A(n914), .B(n915), .Y(n913) );
  OAI221XL U1208 ( .A0(n1120), .A1(n171), .B0(n104), .B1(n18), .C0(n1121), .Y(
        n1583) );
  XNOR2X1 U1209 ( .A(round_key[2]), .B(block[2]), .Y(n1120) );
  AOI222XL U1210 ( .A0(n14), .A1(new_sboxw[2]), .B0(n135), .B1(n459), .C0(n66), 
        .C1(n1122), .Y(n1121) );
  XOR2X1 U1211 ( .A(n1123), .B(n1124), .Y(n1122) );
  OAI221XL U1212 ( .A0(n1303), .A1(n166), .B0(n35), .B1(n10), .C0(n1304), .Y(
        n1601) );
  XNOR2X1 U1213 ( .A(round_key[48]), .B(block[48]), .Y(n1303) );
  AOI222XL U1214 ( .A0(n5), .A1(new_sboxw[16]), .B0(n120), .B1(n774), .C0(n61), 
        .C1(n1305), .Y(n1304) );
  XOR2X1 U1215 ( .A(n1306), .B(n1307), .Y(n1305) );
  OAI221XL U1216 ( .A0(n1138), .A1(n171), .B0(n106), .B1(n18), .C0(n1139), .Y(
        n1585) );
  XNOR2X1 U1217 ( .A(round_key[0]), .B(block[0]), .Y(n1138) );
  AOI222XL U1218 ( .A0(n14), .A1(new_sboxw[0]), .B0(n144), .B1(n1140), .C0(n66), .C1(n1141), .Y(n1139) );
  XOR2X1 U1219 ( .A(n1142), .B(n1143), .Y(n1141) );
  OAI221XL U1220 ( .A0(n1224), .A1(n170), .B0(n24), .B1(n12), .C0(n1225), .Y(
        n1593) );
  XNOR2X1 U1221 ( .A(round_key[24]), .B(block[24]), .Y(n1224) );
  AOI222XL U1222 ( .A0(n6), .A1(new_sboxw[24]), .B0(n116), .B1(n773), .C0(n64), 
        .C1(n1226), .Y(n1225) );
  XOR2X1 U1223 ( .A(n1227), .B(n1228), .Y(n1226) );
  OAI221XL U1224 ( .A0(n983), .A1(n174), .B0(n81), .B1(n19), .C0(n984), .Y(
        n1567) );
  XNOR2X1 U1225 ( .A(round_key[82]), .B(block[82]), .Y(n983) );
  AOI222XL U1226 ( .A0(n15), .A1(new_sboxw[18]), .B0(n147), .B1(n833), .C0(n74), .C1(n985), .Y(n984) );
  XOR2X1 U1227 ( .A(n986), .B(n987), .Y(n985) );
  OAI221XL U1228 ( .A0(n713), .A1(n190), .B0(n134), .B1(n59), .C0(n714), .Y(
        n1539) );
  XNOR2X1 U1229 ( .A(round_key[14]), .B(block[14]), .Y(n713) );
  AOI222XL U1230 ( .A0(n36), .A1(new_sboxw[14]), .B0(n113), .B1(n1667), .C0(
        n78), .C1(n715), .Y(n714) );
  XOR2X1 U1231 ( .A(n716), .B(n717), .Y(n715) );
  OAI221XL U1232 ( .A0(n1332), .A1(n166), .B0(n41), .B1(n10), .C0(n1333), .Y(
        n1605) );
  XNOR2X1 U1233 ( .A(round_key[76]), .B(block[76]), .Y(n1332) );
  AOI222XL U1234 ( .A0(n5), .A1(new_sboxw[12]), .B0(n120), .B1(n1692), .C0(n61), .C1(n1334), .Y(n1333) );
  XOR2X1 U1235 ( .A(n1335), .B(n1336), .Y(n1334) );
  OAI221XL U1236 ( .A0(n738), .A1(n189), .B0(n138), .B1(n59), .C0(n739), .Y(
        n1542) );
  XNOR2X1 U1237 ( .A(round_key[11]), .B(block[11]), .Y(n738) );
  AOI222XL U1238 ( .A0(n36), .A1(new_sboxw[11]), .B0(n113), .B1(n605), .C0(n77), .C1(n740), .Y(n739) );
  XOR2X1 U1239 ( .A(n741), .B(n742), .Y(n740) );
  OAI221XL U1240 ( .A0(n361), .A1(n194), .B0(n175), .B1(n2), .C0(n362), .Y(
        n1503) );
  XNOR2X1 U1241 ( .A(round_key[19]), .B(block[19]), .Y(n361) );
  AOI222XL U1242 ( .A0(new_sboxw[19]), .A1(n155), .B0(n111), .B1(n1659), .C0(
        n85), .C1(n363), .Y(n362) );
  XOR2X1 U1243 ( .A(n364), .B(n365), .Y(n363) );
  OAI221XL U1244 ( .A0(n1282), .A1(n170), .B0(n32), .B1(n10), .C0(n1283), .Y(
        n1599) );
  XNOR2X1 U1245 ( .A(round_key[50]), .B(block[50]), .Y(n1282) );
  AOI222XL U1246 ( .A0(n5), .A1(new_sboxw[18]), .B0(n120), .B1(n1128), .C0(n64), .C1(n1284), .Y(n1283) );
  XOR2X1 U1247 ( .A(n1285), .B(n1286), .Y(n1284) );
  OAI221XL U1248 ( .A0(n1000), .A1(n174), .B0(n84), .B1(n19), .C0(n1001), .Y(
        n1569) );
  XNOR2X1 U1249 ( .A(round_key[80]), .B(block[80]), .Y(n1000) );
  AOI222XL U1250 ( .A0(n15), .A1(new_sboxw[16]), .B0(n107), .B1(n852), .C0(n74), .C1(n1002), .Y(n1001) );
  XOR2X1 U1251 ( .A(n1003), .B(n1004), .Y(n1002) );
  OAI221XL U1252 ( .A0(n795), .A1(n189), .B0(n145), .B1(n40), .C0(n796), .Y(
        n1548) );
  XNOR2X1 U1253 ( .A(round_key[37]), .B(block[37]), .Y(n795) );
  AOI222XL U1254 ( .A0(n30), .A1(new_sboxw[5]), .B0(n113), .B1(n1671), .C0(n77), .C1(n797), .Y(n796) );
  XOR2X1 U1255 ( .A(n798), .B(n799), .Y(n797) );
  OAI221XL U1256 ( .A0(n1292), .A1(n166), .B0(n34), .B1(n10), .C0(n1293), .Y(
        n1600) );
  XNOR2X1 U1257 ( .A(round_key[49]), .B(block[49]), .Y(n1292) );
  AOI222XL U1258 ( .A0(n5), .A1(new_sboxw[17]), .B0(n120), .B1(n1688), .C0(n61), .C1(n1294), .Y(n1293) );
  XOR2X1 U1259 ( .A(n1295), .B(n1296), .Y(n1294) );
  OAI221XL U1260 ( .A0(n1130), .A1(n171), .B0(n105), .B1(n18), .C0(n1131), .Y(
        n1584) );
  XNOR2X1 U1261 ( .A(round_key[1]), .B(block[1]), .Y(n1130) );
  AOI222XL U1262 ( .A0(n14), .A1(new_sboxw[1]), .B0(n135), .B1(n471), .C0(n66), 
        .C1(n1132), .Y(n1131) );
  XOR2X1 U1263 ( .A(n1133), .B(n1134), .Y(n1132) );
  OAI221XL U1264 ( .A0(n721), .A1(n189), .B0(n136), .B1(n59), .C0(n722), .Y(
        n1540) );
  XNOR2X1 U1265 ( .A(round_key[13]), .B(block[13]), .Y(n721) );
  AOI222XL U1266 ( .A0(n561), .A1(new_sboxw[13]), .B0(n113), .B1(n1668), .C0(
        n77), .C1(n723), .Y(n722) );
  XOR2X1 U1267 ( .A(n724), .B(n725), .Y(n723) );
  OAI221XL U1268 ( .A0(n1346), .A1(n166), .B0(n42), .B1(n10), .C0(n1347), .Y(
        n1606) );
  XNOR2X1 U1269 ( .A(round_key[75]), .B(block[75]), .Y(n1346) );
  AOI222XL U1270 ( .A0(n5), .A1(new_sboxw[11]), .B0(n120), .B1(n1113), .C0(n61), .C1(n1348), .Y(n1347) );
  XOR2X1 U1271 ( .A(n1349), .B(n1350), .Y(n1348) );
  OAI221XL U1272 ( .A0(n1158), .A1(n171), .B0(n13), .B1(n1150), .C0(n1159), 
        .Y(n1587) );
  XNOR2X1 U1273 ( .A(round_key[30]), .B(block[30]), .Y(n1158) );
  AOI222XL U1274 ( .A0(n1152), .A1(new_sboxw[30]), .B0(n144), .B1(n1698), .C0(
        n66), .C1(n1160), .Y(n1159) );
  XOR2X1 U1275 ( .A(n1161), .B(n1162), .Y(n1160) );
  OAI221XL U1276 ( .A0(n1270), .A1(n170), .B0(n31), .B1(n12), .C0(n1271), .Y(
        n1598) );
  XNOR2X1 U1277 ( .A(round_key[51]), .B(block[51]), .Y(n1270) );
  AOI222XL U1278 ( .A0(n5), .A1(new_sboxw[19]), .B0(n120), .B1(n1114), .C0(n64), .C1(n1272), .Y(n1271) );
  XOR2X1 U1279 ( .A(n1273), .B(n1274), .Y(n1272) );
  OAI221XL U1280 ( .A0(n1108), .A1(n171), .B0(n103), .B1(n18), .C0(n1109), .Y(
        n1582) );
  XNOR2X1 U1281 ( .A(round_key[3]), .B(block[3]), .Y(n1108) );
  AOI222XL U1282 ( .A0(n14), .A1(new_sboxw[3]), .B0(n144), .B1(n910), .C0(n66), 
        .C1(n1110), .Y(n1109) );
  XOR2X1 U1283 ( .A(n1111), .B(n1112), .Y(n1110) );
  OAI221XL U1284 ( .A0(n1324), .A1(n166), .B0(n39), .B1(n10), .C0(n1325), .Y(
        n1604) );
  XNOR2X1 U1285 ( .A(round_key[77]), .B(block[77]), .Y(n1324) );
  AOI222XL U1286 ( .A0(n5), .A1(new_sboxw[13]), .B0(n120), .B1(n337), .C0(n61), 
        .C1(n1326), .Y(n1325) );
  XOR2X1 U1287 ( .A(n1327), .B(n1328), .Y(n1326) );
  OAI221XL U1288 ( .A0(n729), .A1(n189), .B0(n137), .B1(n59), .C0(n730), .Y(
        n1541) );
  XNOR2X1 U1289 ( .A(round_key[12]), .B(block[12]), .Y(n729) );
  AOI222XL U1290 ( .A0(n36), .A1(new_sboxw[12]), .B0(n113), .B1(n594), .C0(n77), .C1(n731), .Y(n730) );
  XOR2X1 U1291 ( .A(n732), .B(n733), .Y(n731) );
  OAI221XL U1292 ( .A0(n1359), .A1(n166), .B0(n43), .B1(n10), .C0(n1360), .Y(
        n1607) );
  XNOR2X1 U1293 ( .A(round_key[74]), .B(block[74]), .Y(n1359) );
  AOI222XL U1294 ( .A0(n5), .A1(new_sboxw[10]), .B0(n120), .B1(n1126), .C0(n61), .C1(n1361), .Y(n1360) );
  XOR2X1 U1295 ( .A(n1362), .B(n1363), .Y(n1361) );
  OAI221XL U1296 ( .A0(n1190), .A1(n170), .B0(n21), .B1(n12), .C0(n1191), .Y(
        n1590) );
  XNOR2X1 U1297 ( .A(round_key[27]), .B(block[27]), .Y(n1190) );
  AOI222XL U1298 ( .A0(n6), .A1(new_sboxw[27]), .B0(n116), .B1(n748), .C0(n64), 
        .C1(n1192), .Y(n1191) );
  XOR2X1 U1299 ( .A(n1193), .B(n1194), .Y(n1192) );
  OAI221XL U1300 ( .A0(n1204), .A1(n170), .B0(n22), .B1(n12), .C0(n1205), .Y(
        n1591) );
  XNOR2X1 U1301 ( .A(round_key[26]), .B(block[26]), .Y(n1204) );
  AOI222XL U1302 ( .A0(n6), .A1(new_sboxw[26]), .B0(n116), .B1(n756), .C0(n64), 
        .C1(n1206), .Y(n1205) );
  XOR2X1 U1303 ( .A(n1207), .B(n1208), .Y(n1206) );
  OAI221XL U1304 ( .A0(n1215), .A1(n170), .B0(n23), .B1(n12), .C0(n1216), .Y(
        n1592) );
  XNOR2X1 U1305 ( .A(round_key[25]), .B(block[25]), .Y(n1215) );
  AOI222XL U1306 ( .A0(n6), .A1(new_sboxw[25]), .B0(n116), .B1(n1125), .C0(n64), .C1(n1217), .Y(n1216) );
  XOR2X1 U1307 ( .A(n1218), .B(n1219), .Y(n1217) );
  OAI221XL U1308 ( .A0(n1057), .A1(n172), .B0(n94), .B1(n19), .C0(n1058), .Y(
        n1576) );
  XNOR2X1 U1309 ( .A(round_key[105]), .B(block[105]), .Y(n1057) );
  AOI222XL U1310 ( .A0(n14), .A1(new_sboxw[9]), .B0(n242), .B1(n845), .C0(n72), 
        .C1(n1059), .Y(n1058) );
  XOR2X1 U1311 ( .A(n1060), .B(n1061), .Y(n1059) );
  OAI221XL U1312 ( .A0(n492), .A1(n743), .B0(n191), .B1(n160), .C0(n493), .Y(
        n1516) );
  XNOR2X1 U1313 ( .A(round_key[70]), .B(block[70]), .Y(n492) );
  AOI222XL U1314 ( .A0(new_sboxw[6]), .A1(n153), .B0(n135), .B1(n1662), .C0(
        n85), .C1(n494), .Y(n493) );
  XOR2X1 U1315 ( .A(n495), .B(n496), .Y(n494) );
  OAI221XL U1316 ( .A0(n944), .A1(n174), .B0(n73), .B1(n25), .C0(n945), .Y(
        n1563) );
  XNOR2X1 U1317 ( .A(round_key[86]), .B(block[86]), .Y(n944) );
  AOI222XL U1318 ( .A0(n17), .A1(new_sboxw[22]), .B0(n147), .B1(n1674), .C0(
        n74), .C1(n946), .Y(n945) );
  XOR2X1 U1319 ( .A(n947), .B(n948), .Y(n946) );
  OAI221XL U1320 ( .A0(n1400), .A1(n1486), .B0(n48), .B1(n9), .C0(n1401), .Y(
        n1612) );
  XNOR2X1 U1321 ( .A(round_key[101]), .B(block[101]), .Y(n1400) );
  AOI222XL U1322 ( .A0(n4), .A1(new_sboxw[5]), .B0(n128), .B1(n348), .C0(n97), 
        .C1(n1402), .Y(n1401) );
  XOR2X1 U1323 ( .A(n1403), .B(n1404), .Y(n1402) );
  OAI221XL U1324 ( .A0(n1462), .A1(n1486), .B0(n53), .B1(n9), .C0(n1463), .Y(
        n1617) );
  XNOR2X1 U1325 ( .A(round_key[96]), .B(block[96]), .Y(n1462) );
  AOI222XL U1326 ( .A0(n4), .A1(new_sboxw[0]), .B0(n128), .B1(n1201), .C0(n97), 
        .C1(n1464), .Y(n1463) );
  XOR2X1 U1327 ( .A(n1465), .B(n1466), .Y(n1464) );
  OAI221XL U1328 ( .A0(n1441), .A1(n1486), .B0(n51), .B1(n9), .C0(n1442), .Y(
        n1615) );
  XNOR2X1 U1329 ( .A(round_key[98]), .B(block[98]), .Y(n1441) );
  AOI222XL U1330 ( .A0(n4), .A1(new_sboxw[2]), .B0(n128), .B1(n381), .C0(n97), 
        .C1(n1443), .Y(n1442) );
  XOR2X1 U1331 ( .A(n1444), .B(n1445), .Y(n1443) );
  OAI221XL U1332 ( .A0(n1246), .A1(n170), .B0(n28), .B1(n12), .C0(n1247), .Y(
        n1596) );
  XNOR2X1 U1333 ( .A(round_key[53]), .B(block[53]), .Y(n1246) );
  AOI222XL U1334 ( .A0(n6), .A1(new_sboxw[21]), .B0(n116), .B1(n341), .C0(n64), 
        .C1(n1248), .Y(n1247) );
  XOR2X1 U1335 ( .A(n1249), .B(n1250), .Y(n1248) );
  OAI221XL U1336 ( .A0(n1429), .A1(n1486), .B0(n50), .B1(n9), .C0(n1430), .Y(
        n1614) );
  XNOR2X1 U1337 ( .A(round_key[99]), .B(block[99]), .Y(n1429) );
  AOI222XL U1338 ( .A0(n4), .A1(new_sboxw[3]), .B0(n128), .B1(n747), .C0(n97), 
        .C1(n1431), .Y(n1430) );
  XOR2X1 U1339 ( .A(n1432), .B(n1433), .Y(n1431) );
  OAI221XL U1340 ( .A0(n1368), .A1(n166), .B0(n44), .B1(n10), .C0(n1369), .Y(
        n1608) );
  XNOR2X1 U1341 ( .A(round_key[73]), .B(block[73]), .Y(n1368) );
  AOI222XL U1342 ( .A0(n4), .A1(new_sboxw[9]), .B0(n128), .B1(n392), .C0(n61), 
        .C1(n1370), .Y(n1369) );
  XOR2X1 U1343 ( .A(n1371), .B(n1372), .Y(n1370) );
  OAI221XL U1344 ( .A0(n749), .A1(n189), .B0(n139), .B1(n59), .C0(n750), .Y(
        n1543) );
  XNOR2X1 U1345 ( .A(round_key[10]), .B(block[10]), .Y(n749) );
  AOI222XL U1346 ( .A0(n561), .A1(new_sboxw[10]), .B0(n113), .B1(n545), .C0(
        n77), .C1(n751), .Y(n750) );
  XOR2X1 U1347 ( .A(n752), .B(n753), .Y(n751) );
  OAI221XL U1348 ( .A0(n757), .A1(n189), .B0(n140), .B1(n59), .C0(n758), .Y(
        n1544) );
  XNOR2X1 U1349 ( .A(round_key[9]), .B(block[9]), .Y(n757) );
  AOI222XL U1350 ( .A0(n30), .A1(new_sboxw[9]), .B0(n113), .B1(n556), .C0(n77), 
        .C1(n759), .Y(n758) );
  XOR2X1 U1351 ( .A(n760), .B(n761), .Y(n759) );
  OAI221XL U1352 ( .A0(n1166), .A1(n171), .B0(n16), .B1(n1150), .C0(n1167), 
        .Y(n1588) );
  XNOR2X1 U1353 ( .A(round_key[29]), .B(block[29]), .Y(n1166) );
  AOI222XL U1354 ( .A0(n6), .A1(new_sboxw[29]), .B0(n116), .B1(n1699), .C0(n66), .C1(n1168), .Y(n1167) );
  XOR2X1 U1355 ( .A(n1169), .B(n1170), .Y(n1168) );
  OAI221XL U1356 ( .A0(n1470), .A1(n1486), .B0(n199), .B1(n160), .C0(n1471), 
        .Y(n1618) );
  XNOR2X1 U1357 ( .A(round_key[64]), .B(block[64]), .Y(n1470) );
  AOI222XL U1358 ( .A0(new_sboxw[0]), .A1(n153), .B0(n108), .B1(n1071), .C0(
        n97), .C1(n1472), .Y(n1471) );
  XOR2X1 U1359 ( .A(n1004), .B(n1473), .Y(n1472) );
  OAI221XL U1360 ( .A0(n1450), .A1(n1486), .B0(n52), .B1(n9), .C0(n1451), .Y(
        n1616) );
  XNOR2X1 U1361 ( .A(round_key[97]), .B(block[97]), .Y(n1450) );
  AOI222XL U1362 ( .A0(n4), .A1(new_sboxw[1]), .B0(n128), .B1(n755), .C0(n97), 
        .C1(n1452), .Y(n1451) );
  XOR2X1 U1363 ( .A(n1453), .B(n1454), .Y(n1452) );
  XNOR2X1 U1364 ( .A(n123), .B(round_key[86]), .Y(n498) );
  XNOR2X1 U1365 ( .A(n122), .B(round_key[87]), .Y(n637) );
  XNOR2X1 U1366 ( .A(n109), .B(round_key[95]), .Y(n562) );
  XNOR2X1 U1367 ( .A(n71), .B(round_key[55]), .Y(n935) );
  XOR2X1 U1368 ( .A(n16), .B(round_key[29]), .Y(n1086) );
  XOR2X1 U1369 ( .A(n11), .B(round_key[31]), .Y(n1203) );
  XOR2X1 U1370 ( .A(n136), .B(round_key[77]), .Y(n949) );
  XOR2X1 U1371 ( .A(new_block[37]), .B(round_key[37]), .Y(n418) );
  OA22X1 U1372 ( .A0(n1631), .A1(n134), .B0(n205), .B1(n87), .Y(n231) );
  XOR2X1 U1373 ( .A(n145), .B(round_key[69]), .Y(n1322) );
  XOR2X1 U1374 ( .A(n89), .B(round_key[45]), .Y(n1244) );
  XOR2X1 U1375 ( .A(n98), .B(round_key[39]), .Y(n858) );
  XOR2X1 U1376 ( .A(n163), .B(round_key[121]), .Y(n1427) );
  XOR2X1 U1377 ( .A(n20), .B(round_key[28]), .Y(n1163) );
  XOR2X1 U1378 ( .A(new_block[117]), .B(round_key[117]), .Y(n258) );
  XOR2X1 U1379 ( .A(n193), .B(round_key[101]), .Y(n1437) );
  XOR2X1 U1380 ( .A(n129), .B(round_key[81]), .Y(n989) );
  XOR2X1 U1381 ( .A(n73), .B(round_key[54]), .Y(n794) );
  XOR2X1 U1382 ( .A(n191), .B(round_key[102]), .Y(n1420) );
  XOR2X1 U1383 ( .A(n92), .B(round_key[43]), .Y(n1048) );
  XOR2X1 U1384 ( .A(n34), .B(round_key[17]), .Y(n765) );
  XOR2X1 U1385 ( .A(n175), .B(round_key[115]), .Y(n372) );
  XOR2X1 U1386 ( .A(n79), .B(round_key[52]), .Y(n970) );
  XOR2X1 U1387 ( .A(n148), .B(round_key[67]), .Y(n978) );
  XOR2X1 U1388 ( .A(n195), .B(round_key[100]), .Y(n1028) );
  XOR2X1 U1389 ( .A(new_block[70]), .B(round_key[70]), .Y(n788) );
  XOR2X1 U1390 ( .A(n167), .B(round_key[119]), .Y(n1419) );
  XOR2X1 U1391 ( .A(new_block[61]), .B(round_key[61]), .Y(n427) );
  XOR2X1 U1392 ( .A(n121), .B(round_key[88]), .Y(n1005) );
  XOR2X1 U1393 ( .A(new_block[85]), .B(round_key[85]), .Y(n507) );
  XOR2X1 U1394 ( .A(n173), .B(round_key[116]), .Y(n658) );
  XOR2X1 U1395 ( .A(n102), .B(round_key[36]), .Y(n802) );
  XOR2X1 U1396 ( .A(n37), .B(round_key[15]), .Y(n1156) );
  XOR2X1 U1397 ( .A(n41), .B(round_key[12]), .Y(n728) );
  XOR2X1 U1398 ( .A(new_block[93]), .B(round_key[93]), .Y(n497) );
  XOR2X1 U1399 ( .A(new_block[13]), .B(round_key[13]), .Y(n337) );
  XNOR2X1 U1400 ( .A(n137), .B(round_key[76]), .Y(n594) );
  XNOR2X1 U1401 ( .A(n158), .B(round_key[124]), .Y(n270) );
  XNOR2X1 U1402 ( .A(n90), .B(round_key[44]), .Y(n429) );
  XNOR2X1 U1403 ( .A(n94), .B(round_key[41]), .Y(n845) );
  XNOR2X1 U1404 ( .A(n29), .B(round_key[20]), .Y(n350) );
  XNOR2X1 U1405 ( .A(n151), .B(round_key[64]), .Y(n633) );
  XOR2X1 U1406 ( .A(new_block[16]), .B(round_key[16]), .Y(n774) );
  XNOR2X1 U1407 ( .A(n146), .B(round_key[68]), .Y(n509) );
  XOR2X1 U1408 ( .A(new_block[92]), .B(round_key[92]), .Y(n510) );
  XOR2X1 U1409 ( .A(new_block[120]), .B(round_key[120]), .Y(n314) );
  XNOR2X1 U1410 ( .A(n105), .B(round_key[33]), .Y(n471) );
  XNOR2X1 U1411 ( .A(n198), .B(round_key[97]), .Y(n310) );
  XNOR2X1 U1412 ( .A(n150), .B(round_key[65]), .Y(n546) );
  XNOR2X1 U1413 ( .A(n28), .B(round_key[21]), .Y(n341) );
  XNOR2X1 U1414 ( .A(n44), .B(round_key[9]), .Y(n392) );
  XOR2X1 U1415 ( .A(new_block[109]), .B(round_key[109]), .Y(n268) );
  XOR2X1 U1416 ( .A(new_block[5]), .B(round_key[5]), .Y(n348) );
  XOR2X1 U1417 ( .A(new_block[1]), .B(round_key[1]), .Y(n755) );
  XOR2X1 U1418 ( .A(new_block[105]), .B(round_key[105]), .Y(n463) );
  XOR2X1 U1419 ( .A(new_block[73]), .B(round_key[73]), .Y(n556) );
  XNOR2X1 U1420 ( .A(n23), .B(round_key[25]), .Y(n1125) );
  XOR2X1 U1421 ( .A(new_block[60]), .B(round_key[60]), .Y(n439) );
  XOR2X1 U1422 ( .A(new_block[125]), .B(round_key[125]), .Y(n261) );
  XOR2X1 U1423 ( .A(new_block[89]), .B(round_key[89]), .Y(n543) );
  XOR2X1 U1424 ( .A(new_block[57]), .B(round_key[57]), .Y(n834) );
  XOR2X1 U1425 ( .A(new_block[108]), .B(round_key[108]), .Y(n280) );
  XOR2X1 U1426 ( .A(new_block[4]), .B(round_key[4]), .Y(n360) );
  XOR2X1 U1427 ( .A(new_block[84]), .B(round_key[84]), .Y(n520) );
  XOR2X1 U1428 ( .A(new_block[113]), .B(round_key[113]), .Y(n300) );
  XNOR2X1 U1429 ( .A(n161), .B(round_key[122]), .Y(n294) );
  XNOR2X1 U1430 ( .A(n67), .B(round_key[59]), .Y(n821) );
  XOR2X1 U1431 ( .A(new_block[56]), .B(round_key[56]), .Y(n853) );
  XOR2X1 U1432 ( .A(new_block[91]), .B(round_key[91]), .Y(n597) );
  XOR2X1 U1433 ( .A(new_block[27]), .B(round_key[27]), .Y(n748) );
  XOR2X1 U1434 ( .A(new_block[26]), .B(round_key[26]), .Y(n756) );
  XNOR2X1 U1435 ( .A(n185), .B(round_key[106]), .Y(n452) );
  XNOR2X1 U1436 ( .A(n68), .B(round_key[58]), .Y(n832) );
  XNOR2X1 U1437 ( .A(n159), .B(round_key[123]), .Y(n283) );
  XOR2X1 U1438 ( .A(new_block[90]), .B(round_key[90]), .Y(n609) );
  XNOR2X1 U1439 ( .A(n43), .B(round_key[10]), .Y(n1126) );
  XOR2X1 U1440 ( .A(new_block[51]), .B(round_key[51]), .Y(n822) );
  XNOR2X1 U1441 ( .A(n126), .B(round_key[83]), .Y(n604) );
  XNOR2X1 U1442 ( .A(n93), .B(round_key[42]), .Y(n836) );
  XNOR2X1 U1443 ( .A(n149), .B(round_key[66]), .Y(n825) );
  XNOR2X1 U1444 ( .A(n84), .B(round_key[48]), .Y(n852) );
  XOR2X1 U1445 ( .A(new_block[98]), .B(round_key[98]), .Y(n535) );
  XOR2X1 U1446 ( .A(new_block[104]), .B(round_key[104]), .Y(n475) );
  XOR2X1 U1447 ( .A(new_block[2]), .B(round_key[2]), .Y(n381) );
  XOR2X1 U1448 ( .A(new_block[50]), .B(round_key[50]), .Y(n833) );
  XNOR2X1 U1449 ( .A(n50), .B(round_key[3]), .Y(n747) );
  XOR2X1 U1450 ( .A(new_block[99]), .B(round_key[99]), .Y(n523) );
  XOR2X1 U1451 ( .A(new_block[74]), .B(round_key[74]), .Y(n545) );
  XOR2X1 U1452 ( .A(new_block[40]), .B(round_key[40]), .Y(n854) );
  XOR2X1 U1453 ( .A(new_block[34]), .B(round_key[34]), .Y(n459) );
  XOR2X1 U1454 ( .A(new_block[24]), .B(round_key[24]), .Y(n773) );
  XOR2X1 U1455 ( .A(new_block[82]), .B(round_key[82]), .Y(n616) );
  XOR2X1 U1456 ( .A(new_block[8]), .B(round_key[8]), .Y(n1147) );
  XOR2X1 U1457 ( .A(new_block[114]), .B(round_key[114]), .Y(n302) );
  XOR2X1 U1458 ( .A(new_block[112]), .B(round_key[112]), .Y(n396) );
  XOR2X1 U1459 ( .A(new_block[18]), .B(round_key[18]), .Y(n1128) );
  XNOR2X1 U1460 ( .A(n53), .B(round_key[0]), .Y(n1201) );
  XOR2X1 U1461 ( .A(new_block[96]), .B(round_key[96]), .Y(n1071) );
  XOR2X1 U1462 ( .A(new_block[72]), .B(round_key[72]), .Y(n768) );
  XOR2X1 U1463 ( .A(new_block[80]), .B(round_key[80]), .Y(n697) );
  XOR2X1 U1464 ( .A(new_block[32]), .B(round_key[32]), .Y(n1140) );
  NOR2X1 U1465 ( .A(n57), .B(sword_ctr_reg[1]), .Y(n862) );
  NOR2X1 U1466 ( .A(n56), .B(n57), .Y(n1469) );
  NOR2X1 U1467 ( .A(n56), .B(sword_ctr_reg[0]), .Y(n1148) );
  OAI221XL U1468 ( .A0(n1638), .A1(n48), .B0(n1636), .B1(n193), .C0(n209), .Y(
        tmp_sboxw[5]) );
  OA22X1 U1469 ( .A0(n1633), .A1(n145), .B0(n1629), .B1(n100), .Y(n209) );
  OAI221XL U1470 ( .A0(n1638), .A1(n16), .B0(n1636), .B1(n157), .C0(n215), .Y(
        tmp_sboxw[29]) );
  OA22X1 U1471 ( .A0(n1633), .A1(n112), .B0(n1629), .B1(n63), .Y(n215) );
  OAI221XL U1472 ( .A0(n201), .A1(n28), .B0(n1635), .B1(n169), .C0(n223), .Y(
        tmp_sboxw[21]) );
  OA22X1 U1473 ( .A0(n1632), .A1(n124), .B0(n1628), .B1(n76), .Y(n223) );
  OAI221XL U1474 ( .A0(n1637), .A1(n39), .B0(n1634), .B1(n182), .C0(n232), .Y(
        tmp_sboxw[13]) );
  OA22X1 U1475 ( .A0(n1631), .A1(n136), .B0(n205), .B1(n89), .Y(n232) );
  OAI221XL U1476 ( .A0(n237), .A1(n192), .B0(n152), .B1(n2), .C0(n240), .Y(
        n1491) );
  XNOR2X1 U1477 ( .A(round_key[127]), .B(block[127]), .Y(n237) );
  AOI222XL U1478 ( .A0(new_sboxw[31]), .A1(n241), .B0(n115), .B1(n243), .C0(
        n82), .C1(n245), .Y(n240) );
  XOR2X1 U1479 ( .A(n246), .B(n247), .Y(n245) );
  OAI221XL U1480 ( .A0(n271), .A1(n192), .B0(n158), .B1(n165), .C0(n272), .Y(
        n1494) );
  XNOR2X1 U1481 ( .A(round_key[124]), .B(block[124]), .Y(n271) );
  AOI222XL U1482 ( .A0(new_sboxw[28]), .A1(n156), .B0(n108), .B1(n270), .C0(
        n82), .C1(n273), .Y(n272) );
  XOR2X1 U1483 ( .A(n274), .B(n275), .Y(n273) );
  OAI221XL U1484 ( .A0(n322), .A1(n192), .B0(n167), .B1(n165), .C0(n323), .Y(
        n1499) );
  XNOR2X1 U1485 ( .A(round_key[23]), .B(block[23]), .Y(n322) );
  AOI222XL U1486 ( .A0(new_sboxw[23]), .A1(n156), .B0(n111), .B1(n1655), .C0(
        n82), .C1(n324), .Y(n323) );
  XOR2X1 U1487 ( .A(n325), .B(n326), .Y(n324) );
  OAI221XL U1488 ( .A0(n635), .A1(n190), .B0(n122), .B1(n60), .C0(n636), .Y(
        n1530) );
  XNOR2X1 U1489 ( .A(round_key[119]), .B(block[119]), .Y(n635) );
  AOI222XL U1490 ( .A0(n33), .A1(new_sboxw[23]), .B0(n131), .B1(n637), .C0(n78), .C1(n638), .Y(n636) );
  XOR2X1 U1491 ( .A(n639), .B(n640), .Y(n638) );
  OAI221XL U1492 ( .A0(n482), .A1(n194), .B0(n188), .B1(n160), .C0(n483), .Y(
        n1515) );
  XNOR2X1 U1493 ( .A(round_key[71]), .B(block[71]), .Y(n482) );
  AOI222XL U1494 ( .A0(new_sboxw[7]), .A1(n153), .B0(n135), .B1(n484), .C0(n88), .C1(n485), .Y(n483) );
  XOR2X1 U1495 ( .A(n486), .B(n487), .Y(n485) );
  OAI221XL U1496 ( .A0(n558), .A1(n200), .B0(n109), .B1(n559), .C0(n560), .Y(
        n1522) );
  XNOR2X1 U1497 ( .A(round_key[95]), .B(block[95]), .Y(n558) );
  AOI222XL U1498 ( .A0(n36), .A1(new_sboxw[31]), .B0(n131), .B1(n562), .C0(n91), .C1(n563), .Y(n560) );
  XOR2X1 U1499 ( .A(n564), .B(n565), .Y(n563) );
  OAI221XL U1500 ( .A0(n778), .A1(n189), .B0(n142), .B1(n40), .C0(n779), .Y(
        n1546) );
  XNOR2X1 U1501 ( .A(round_key[39]), .B(block[39]), .Y(n778) );
  AOI222XL U1502 ( .A0(n30), .A1(new_sboxw[7]), .B0(n113), .B1(n567), .C0(n77), 
        .C1(n780), .Y(n779) );
  XOR2X1 U1503 ( .A(n781), .B(n782), .Y(n780) );
  OAI221XL U1504 ( .A0(n936), .A1(n174), .B0(n71), .B1(n25), .C0(n937), .Y(
        n1562) );
  XNOR2X1 U1505 ( .A(round_key[87]), .B(block[87]), .Y(n936) );
  AOI222XL U1506 ( .A0(n17), .A1(new_sboxw[23]), .B0(n135), .B1(n935), .C0(n74), .C1(n938), .Y(n937) );
  XOR2X1 U1507 ( .A(n939), .B(n940), .Y(n938) );
  OAI221XL U1508 ( .A0(n1074), .A1(n172), .B0(n98), .B1(n18), .C0(n1075), .Y(
        n1578) );
  XNOR2X1 U1509 ( .A(round_key[7]), .B(block[7]), .Y(n1074) );
  AOI222XL U1510 ( .A0(n14), .A1(new_sboxw[7]), .B0(n144), .B1(n1685), .C0(n72), .C1(n1076), .Y(n1075) );
  XOR2X1 U1511 ( .A(n1077), .B(n1078), .Y(n1076) );
  OAI221XL U1512 ( .A0(n863), .A1(n180), .B0(n58), .B1(n864), .C0(n865), .Y(
        n1554) );
  XNOR2X1 U1513 ( .A(round_key[63]), .B(block[63]), .Y(n863) );
  AOI222XL U1514 ( .A0(n866), .A1(new_sboxw[31]), .B0(n115), .B1(n859), .C0(
        n75), .C1(n867), .Y(n865) );
  XOR2X1 U1515 ( .A(n868), .B(n869), .Y(n867) );
  OAI221XL U1516 ( .A0(n1231), .A1(n170), .B0(n26), .B1(n12), .C0(n1232), .Y(
        n1594) );
  XNOR2X1 U1517 ( .A(round_key[55]), .B(block[55]), .Y(n1231) );
  AOI222XL U1518 ( .A0(n6), .A1(new_sboxw[23]), .B0(n116), .B1(n710), .C0(n64), 
        .C1(n1233), .Y(n1232) );
  XOR2X1 U1519 ( .A(n1234), .B(n1235), .Y(n1233) );
  OAI221XL U1520 ( .A0(n1149), .A1(n171), .B0(n11), .B1(n1150), .C0(n1151), 
        .Y(n1586) );
  XNOR2X1 U1521 ( .A(round_key[31]), .B(block[31]), .Y(n1149) );
  AOI222XL U1522 ( .A0(n1152), .A1(new_sboxw[31]), .B0(n107), .B1(n1694), .C0(
        n66), .C1(n1153), .Y(n1151) );
  XOR2X1 U1523 ( .A(n1154), .B(n1155), .Y(n1153) );
  OAI221XL U1524 ( .A0(n1387), .A1(n1486), .B0(n46), .B1(n9), .C0(n1388), .Y(
        n1610) );
  XNOR2X1 U1525 ( .A(round_key[103]), .B(block[103]), .Y(n1387) );
  AOI222XL U1526 ( .A0(n4), .A1(new_sboxw[7]), .B0(n128), .B1(n777), .C0(n97), 
        .C1(n1389), .Y(n1388) );
  XOR2X1 U1527 ( .A(n1390), .B(n1011), .Y(n1389) );
  OAI221XL U1528 ( .A0(n659), .A1(n190), .B0(n125), .B1(n60), .C0(n660), .Y(
        n1533) );
  XNOR2X1 U1529 ( .A(round_key[116]), .B(block[116]), .Y(n659) );
  AOI222XL U1530 ( .A0(n33), .A1(new_sboxw[20]), .B0(n144), .B1(n520), .C0(n78), .C1(n661), .Y(n660) );
  XOR2X1 U1531 ( .A(n662), .B(n663), .Y(n661) );
  OAI221XL U1532 ( .A0(n960), .A1(n174), .B0(n79), .B1(n25), .C0(n961), .Y(
        n1565) );
  XNOR2X1 U1533 ( .A(round_key[84]), .B(block[84]), .Y(n960) );
  AOI222XL U1534 ( .A0(n17), .A1(new_sboxw[20]), .B0(n147), .B1(n1678), .C0(
        n74), .C1(n962), .Y(n961) );
  XOR2X1 U1535 ( .A(n963), .B(n964), .Y(n962) );
  OAI221XL U1536 ( .A0(n511), .A1(n200), .B0(n195), .B1(n160), .C0(n512), .Y(
        n1518) );
  XNOR2X1 U1537 ( .A(round_key[68]), .B(block[68]), .Y(n511) );
  AOI222XL U1538 ( .A0(new_sboxw[4]), .A1(n153), .B0(n101), .B1(n1664), .C0(
        n91), .C1(n513), .Y(n512) );
  XOR2X1 U1539 ( .A(n514), .B(n515), .Y(n513) );
  OAI221XL U1540 ( .A0(n585), .A1(n200), .B0(n114), .B1(n60), .C0(n586), .Y(
        n1525) );
  XNOR2X1 U1541 ( .A(round_key[92]), .B(block[92]), .Y(n585) );
  AOI222XL U1542 ( .A0(n33), .A1(new_sboxw[28]), .B0(n131), .B1(n510), .C0(n85), .C1(n587), .Y(n586) );
  XOR2X1 U1543 ( .A(n588), .B(n589), .Y(n587) );
  OAI221XL U1544 ( .A0(n803), .A1(n189), .B0(n146), .B1(n40), .C0(n804), .Y(
        n1549) );
  XNOR2X1 U1545 ( .A(round_key[36]), .B(block[36]), .Y(n803) );
  AOI222XL U1546 ( .A0(n30), .A1(new_sboxw[4]), .B0(n115), .B1(n509), .C0(n77), 
        .C1(n805), .Y(n804) );
  XOR2X1 U1547 ( .A(n806), .B(n807), .Y(n805) );
  OAI221XL U1548 ( .A0(n889), .A1(n180), .B0(n65), .B1(n25), .C0(n890), .Y(
        n1557) );
  XNOR2X1 U1549 ( .A(round_key[60]), .B(block[60]), .Y(n889) );
  AOI222XL U1550 ( .A0(n17), .A1(new_sboxw[28]), .B0(n115), .B1(n439), .C0(n75), .C1(n891), .Y(n890) );
  XOR2X1 U1551 ( .A(n892), .B(n893), .Y(n891) );
  OAI221XL U1552 ( .A0(n351), .A1(n239), .B0(n173), .B1(n165), .C0(n352), .Y(
        n1502) );
  XNOR2X1 U1553 ( .A(round_key[20]), .B(block[20]), .Y(n351) );
  AOI222XL U1554 ( .A0(new_sboxw[20]), .A1(n156), .B0(n111), .B1(n1658), .C0(
        n85), .C1(n353), .Y(n352) );
  XOR2X1 U1555 ( .A(n354), .B(n355), .Y(n353) );
  OAI221XL U1556 ( .A0(n1411), .A1(n1486), .B0(n49), .B1(n9), .C0(n1412), .Y(
        n1613) );
  XNOR2X1 U1557 ( .A(round_key[100]), .B(block[100]), .Y(n1411) );
  AOI222XL U1558 ( .A0(n4), .A1(new_sboxw[4]), .B0(n128), .B1(n360), .C0(n97), 
        .C1(n1413), .Y(n1412) );
  XOR2X1 U1559 ( .A(n1414), .B(n1415), .Y(n1413) );
  OAI221XL U1560 ( .A0(n1256), .A1(n170), .B0(n29), .B1(n12), .C0(n1257), .Y(
        n1597) );
  XNOR2X1 U1561 ( .A(round_key[52]), .B(block[52]), .Y(n1256) );
  AOI222XL U1562 ( .A0(n6), .A1(new_sboxw[20]), .B0(n116), .B1(n350), .C0(n64), 
        .C1(n1258), .Y(n1257) );
  XOR2X1 U1563 ( .A(n1259), .B(n1260), .Y(n1258) );
  OAI221XL U1564 ( .A0(n1098), .A1(n171), .B0(n102), .B1(n18), .C0(n1099), .Y(
        n1581) );
  XNOR2X1 U1565 ( .A(round_key[4]), .B(block[4]), .Y(n1098) );
  AOI222XL U1566 ( .A0(n14), .A1(new_sboxw[4]), .B0(n242), .B1(n1686), .C0(n66), .C1(n1100), .Y(n1099) );
  XOR2X1 U1567 ( .A(n1101), .B(n1102), .Y(n1100) );
  OAI221XL U1568 ( .A0(n1176), .A1(n171), .B0(n20), .B1(n12), .C0(n1177), .Y(
        n1589) );
  XNOR2X1 U1569 ( .A(round_key[28]), .B(block[28]), .Y(n1176) );
  AOI222XL U1570 ( .A0(n6), .A1(new_sboxw[28]), .B0(n116), .B1(n1700), .C0(n66), .C1(n1178), .Y(n1177) );
  XOR2X1 U1571 ( .A(n1179), .B(n1180), .Y(n1178) );
  XOR2X1 U1572 ( .A(new_block[107]), .B(round_key[107]), .Y(n442) );
  XOR2X1 U1573 ( .A(new_block[11]), .B(round_key[11]), .Y(n1113) );
  XOR2X1 U1574 ( .A(new_block[35]), .B(round_key[35]), .Y(n910) );
  XOR2X1 U1575 ( .A(new_block[75]), .B(round_key[75]), .Y(n605) );
  XOR2X1 U1576 ( .A(new_block[19]), .B(round_key[19]), .Y(n1114) );
  OA22X1 U1577 ( .A0(n1631), .A1(n132), .B0(n1630), .B1(n86), .Y(n230) );
  OAI221XL U1578 ( .A0(n201), .A1(n27), .B0(n1635), .B1(n168), .C0(n222), .Y(
        tmp_sboxw[22]) );
  OA22X1 U1579 ( .A0(n1632), .A1(n123), .B0(n1628), .B1(n73), .Y(n222) );
  OAI221XL U1580 ( .A0(n1638), .A1(n13), .B0(n1636), .B1(n154), .C0(n213), .Y(
        tmp_sboxw[30]) );
  OA22X1 U1581 ( .A0(n1633), .A1(n110), .B0(n1629), .B1(n62), .Y(n213) );
  OAI221XL U1582 ( .A0(n201), .A1(n26), .B0(n1635), .B1(n167), .C0(n221), .Y(
        tmp_sboxw[23]) );
  OA22X1 U1583 ( .A0(n1632), .A1(n122), .B0(n1628), .B1(n71), .Y(n221) );
  OAI221XL U1584 ( .A0(n1638), .A1(n11), .B0(n1636), .B1(n152), .C0(n212), .Y(
        tmp_sboxw[31]) );
  OA22X1 U1585 ( .A0(n1633), .A1(n109), .B0(n1629), .B1(n58), .Y(n212) );
  OAI221XL U1586 ( .A0(n1638), .A1(n47), .B0(n1636), .B1(n191), .C0(n208), .Y(
        tmp_sboxw[6]) );
  OA22X1 U1587 ( .A0(n1633), .A1(n143), .B0(n1629), .B1(n99), .Y(n208) );
  OAI221XL U1588 ( .A0(n1639), .A1(n46), .B0(n202), .B1(n188), .C0(n207), .Y(
        tmp_sboxw[7]) );
  OA22X1 U1589 ( .A0(n204), .A1(n142), .B0(n1630), .B1(n98), .Y(n207) );
  OAI22XL U1590 ( .A0(n56), .A1(n1487), .B0(n1488), .B1(n1706), .Y(n1626) );
  NOR2X1 U1591 ( .A(n862), .B(n1148), .Y(n1488) );
  OAI22XL U1592 ( .A0(n57), .A1(n1487), .B0(sword_ctr_reg[0]), .B1(n1706), .Y(
        n1627) );
  OAI21XL U1593 ( .A0(n1483), .A1(n54), .B0(n1484), .Y(n1480) );
  NAND3X1 U1594 ( .A(n8), .B(n7), .C(next), .Y(n1478) );
  AOI2BB1X1 U1595 ( .A0N(n1483), .A1N(n55), .B0(n1703), .Y(n1484) );
  OAI21XL U1596 ( .A0(n55), .A1(n1485), .B0(n1482), .Y(n1623) );
  NAND2X1 U1597 ( .A(n8), .B(n1706), .Y(n1487) );
  OR2X1 U1598 ( .A(n1483), .B(round[0]), .Y(n1482) );
  AO21X1 U1599 ( .A0(n1480), .A1(round[2]), .B0(n1481), .Y(n1621) );
  OAI32X1 U1600 ( .A0(round[1]), .A1(round[2]), .A2(n1482), .B0(n1708), .B1(
        n1478), .Y(n1481) );
  INVXL U1601 ( .A(keylen), .Y(n1708) );
  AO21X1 U1602 ( .A0(ready), .A1(n1478), .B0(n108), .Y(n1619) );
  OAI221XL U1603 ( .A0(round[1]), .A1(n1482), .B0(n1484), .B1(n54), .C0(n1478), 
        .Y(n1622) );
  OAI211X1 U1604 ( .A0(n1702), .A1(n7), .B0(n1475), .C0(n1483), .Y(n1625) );
  OAI211X1 U1605 ( .A0(n1703), .A1(n1476), .B0(n1478), .C0(n1479), .Y(n1620)
         );
  OAI21XL U1606 ( .A0(round[2]), .A1(n1480), .B0(round[3]), .Y(n1479) );
  OAI211X1 U1607 ( .A0(n1702), .A1(n8), .B0(n1483), .C0(n1478), .Y(n1624) );
  INVX1 U1608 ( .A(n1490), .Y(n1702) );
  AOI221XL U1609 ( .A0(n1489), .A1(n1469), .B0(n7), .B1(next), .C0(
        \dec_ctrl_reg[0] ), .Y(n1490) );
endmodule


module aes_key_mem ( clk, reset_n, key, keylen, init, round, round_key, ready, 
        sboxw, new_sboxw );
  input [255:0] key;
  input [3:0] round;
  output [127:0] round_key;
  output [31:0] sboxw;
  input [31:0] new_sboxw;
  input clk, reset_n, keylen, init;
  output ready;
  wire   N31, N32, N33, N34, \key_mem[0][127] , \key_mem[0][126] ,
         \key_mem[0][125] , \key_mem[0][124] , \key_mem[0][123] ,
         \key_mem[0][122] , \key_mem[0][121] , \key_mem[0][120] ,
         \key_mem[0][119] , \key_mem[0][118] , \key_mem[0][117] ,
         \key_mem[0][116] , \key_mem[0][115] , \key_mem[0][114] ,
         \key_mem[0][113] , \key_mem[0][112] , \key_mem[0][111] ,
         \key_mem[0][110] , \key_mem[0][109] , \key_mem[0][108] ,
         \key_mem[0][107] , \key_mem[0][106] , \key_mem[0][105] ,
         \key_mem[0][104] , \key_mem[0][103] , \key_mem[0][102] ,
         \key_mem[0][101] , \key_mem[0][100] , \key_mem[0][99] ,
         \key_mem[0][98] , \key_mem[0][97] , \key_mem[0][96] ,
         \key_mem[0][95] , \key_mem[0][94] , \key_mem[0][93] ,
         \key_mem[0][92] , \key_mem[0][91] , \key_mem[0][90] ,
         \key_mem[0][89] , \key_mem[0][88] , \key_mem[0][87] ,
         \key_mem[0][86] , \key_mem[0][85] , \key_mem[0][84] ,
         \key_mem[0][83] , \key_mem[0][82] , \key_mem[0][81] ,
         \key_mem[0][80] , \key_mem[0][79] , \key_mem[0][78] ,
         \key_mem[0][77] , \key_mem[0][76] , \key_mem[0][75] ,
         \key_mem[0][74] , \key_mem[0][73] , \key_mem[0][72] ,
         \key_mem[0][71] , \key_mem[0][70] , \key_mem[0][69] ,
         \key_mem[0][68] , \key_mem[0][67] , \key_mem[0][66] ,
         \key_mem[0][65] , \key_mem[0][64] , \key_mem[0][63] ,
         \key_mem[0][62] , \key_mem[0][61] , \key_mem[0][60] ,
         \key_mem[0][59] , \key_mem[0][58] , \key_mem[0][57] ,
         \key_mem[0][56] , \key_mem[0][55] , \key_mem[0][54] ,
         \key_mem[0][53] , \key_mem[0][52] , \key_mem[0][51] ,
         \key_mem[0][50] , \key_mem[0][49] , \key_mem[0][48] ,
         \key_mem[0][47] , \key_mem[0][46] , \key_mem[0][45] ,
         \key_mem[0][44] , \key_mem[0][43] , \key_mem[0][42] ,
         \key_mem[0][41] , \key_mem[0][40] , \key_mem[0][39] ,
         \key_mem[0][38] , \key_mem[0][37] , \key_mem[0][36] ,
         \key_mem[0][35] , \key_mem[0][34] , \key_mem[0][33] ,
         \key_mem[0][32] , \key_mem[0][31] , \key_mem[0][30] ,
         \key_mem[0][29] , \key_mem[0][28] , \key_mem[0][27] ,
         \key_mem[0][26] , \key_mem[0][25] , \key_mem[0][24] ,
         \key_mem[0][23] , \key_mem[0][22] , \key_mem[0][21] ,
         \key_mem[0][20] , \key_mem[0][19] , \key_mem[0][18] ,
         \key_mem[0][17] , \key_mem[0][16] , \key_mem[0][15] ,
         \key_mem[0][14] , \key_mem[0][13] , \key_mem[0][12] ,
         \key_mem[0][11] , \key_mem[0][10] , \key_mem[0][9] , \key_mem[0][8] ,
         \key_mem[0][7] , \key_mem[0][6] , \key_mem[0][5] , \key_mem[0][4] ,
         \key_mem[0][3] , \key_mem[0][2] , \key_mem[0][1] , \key_mem[0][0] ,
         \key_mem[1][127] , \key_mem[1][126] , \key_mem[1][125] ,
         \key_mem[1][124] , \key_mem[1][123] , \key_mem[1][122] ,
         \key_mem[1][121] , \key_mem[1][120] , \key_mem[1][119] ,
         \key_mem[1][118] , \key_mem[1][117] , \key_mem[1][116] ,
         \key_mem[1][115] , \key_mem[1][114] , \key_mem[1][113] ,
         \key_mem[1][112] , \key_mem[1][111] , \key_mem[1][110] ,
         \key_mem[1][109] , \key_mem[1][108] , \key_mem[1][107] ,
         \key_mem[1][106] , \key_mem[1][105] , \key_mem[1][104] ,
         \key_mem[1][103] , \key_mem[1][102] , \key_mem[1][101] ,
         \key_mem[1][100] , \key_mem[1][99] , \key_mem[1][98] ,
         \key_mem[1][97] , \key_mem[1][96] , \key_mem[1][95] ,
         \key_mem[1][94] , \key_mem[1][93] , \key_mem[1][92] ,
         \key_mem[1][91] , \key_mem[1][90] , \key_mem[1][89] ,
         \key_mem[1][88] , \key_mem[1][87] , \key_mem[1][86] ,
         \key_mem[1][85] , \key_mem[1][84] , \key_mem[1][83] ,
         \key_mem[1][82] , \key_mem[1][81] , \key_mem[1][80] ,
         \key_mem[1][79] , \key_mem[1][78] , \key_mem[1][77] ,
         \key_mem[1][76] , \key_mem[1][75] , \key_mem[1][74] ,
         \key_mem[1][73] , \key_mem[1][72] , \key_mem[1][71] ,
         \key_mem[1][70] , \key_mem[1][69] , \key_mem[1][68] ,
         \key_mem[1][67] , \key_mem[1][66] , \key_mem[1][65] ,
         \key_mem[1][64] , \key_mem[1][63] , \key_mem[1][62] ,
         \key_mem[1][61] , \key_mem[1][60] , \key_mem[1][59] ,
         \key_mem[1][58] , \key_mem[1][57] , \key_mem[1][56] ,
         \key_mem[1][55] , \key_mem[1][54] , \key_mem[1][53] ,
         \key_mem[1][52] , \key_mem[1][51] , \key_mem[1][50] ,
         \key_mem[1][49] , \key_mem[1][48] , \key_mem[1][47] ,
         \key_mem[1][46] , \key_mem[1][45] , \key_mem[1][44] ,
         \key_mem[1][43] , \key_mem[1][42] , \key_mem[1][41] ,
         \key_mem[1][40] , \key_mem[1][39] , \key_mem[1][38] ,
         \key_mem[1][37] , \key_mem[1][36] , \key_mem[1][35] ,
         \key_mem[1][34] , \key_mem[1][33] , \key_mem[1][32] ,
         \key_mem[1][31] , \key_mem[1][30] , \key_mem[1][29] ,
         \key_mem[1][28] , \key_mem[1][27] , \key_mem[1][26] ,
         \key_mem[1][25] , \key_mem[1][24] , \key_mem[1][23] ,
         \key_mem[1][22] , \key_mem[1][21] , \key_mem[1][20] ,
         \key_mem[1][19] , \key_mem[1][18] , \key_mem[1][17] ,
         \key_mem[1][16] , \key_mem[1][15] , \key_mem[1][14] ,
         \key_mem[1][13] , \key_mem[1][12] , \key_mem[1][11] ,
         \key_mem[1][10] , \key_mem[1][9] , \key_mem[1][8] , \key_mem[1][7] ,
         \key_mem[1][6] , \key_mem[1][5] , \key_mem[1][4] , \key_mem[1][3] ,
         \key_mem[1][2] , \key_mem[1][1] , \key_mem[1][0] , \key_mem[2][127] ,
         \key_mem[2][126] , \key_mem[2][125] , \key_mem[2][124] ,
         \key_mem[2][123] , \key_mem[2][122] , \key_mem[2][121] ,
         \key_mem[2][120] , \key_mem[2][119] , \key_mem[2][118] ,
         \key_mem[2][117] , \key_mem[2][116] , \key_mem[2][115] ,
         \key_mem[2][114] , \key_mem[2][113] , \key_mem[2][112] ,
         \key_mem[2][111] , \key_mem[2][110] , \key_mem[2][109] ,
         \key_mem[2][108] , \key_mem[2][107] , \key_mem[2][106] ,
         \key_mem[2][105] , \key_mem[2][104] , \key_mem[2][103] ,
         \key_mem[2][102] , \key_mem[2][101] , \key_mem[2][100] ,
         \key_mem[2][99] , \key_mem[2][98] , \key_mem[2][97] ,
         \key_mem[2][96] , \key_mem[2][95] , \key_mem[2][94] ,
         \key_mem[2][93] , \key_mem[2][92] , \key_mem[2][91] ,
         \key_mem[2][90] , \key_mem[2][89] , \key_mem[2][88] ,
         \key_mem[2][87] , \key_mem[2][86] , \key_mem[2][85] ,
         \key_mem[2][84] , \key_mem[2][83] , \key_mem[2][82] ,
         \key_mem[2][81] , \key_mem[2][80] , \key_mem[2][79] ,
         \key_mem[2][78] , \key_mem[2][77] , \key_mem[2][76] ,
         \key_mem[2][75] , \key_mem[2][74] , \key_mem[2][73] ,
         \key_mem[2][72] , \key_mem[2][71] , \key_mem[2][70] ,
         \key_mem[2][69] , \key_mem[2][68] , \key_mem[2][67] ,
         \key_mem[2][66] , \key_mem[2][65] , \key_mem[2][64] ,
         \key_mem[2][63] , \key_mem[2][62] , \key_mem[2][61] ,
         \key_mem[2][60] , \key_mem[2][59] , \key_mem[2][58] ,
         \key_mem[2][57] , \key_mem[2][56] , \key_mem[2][55] ,
         \key_mem[2][54] , \key_mem[2][53] , \key_mem[2][52] ,
         \key_mem[2][51] , \key_mem[2][50] , \key_mem[2][49] ,
         \key_mem[2][48] , \key_mem[2][47] , \key_mem[2][46] ,
         \key_mem[2][45] , \key_mem[2][44] , \key_mem[2][43] ,
         \key_mem[2][42] , \key_mem[2][41] , \key_mem[2][40] ,
         \key_mem[2][39] , \key_mem[2][38] , \key_mem[2][37] ,
         \key_mem[2][36] , \key_mem[2][35] , \key_mem[2][34] ,
         \key_mem[2][33] , \key_mem[2][32] , \key_mem[2][31] ,
         \key_mem[2][30] , \key_mem[2][29] , \key_mem[2][28] ,
         \key_mem[2][27] , \key_mem[2][26] , \key_mem[2][25] ,
         \key_mem[2][24] , \key_mem[2][23] , \key_mem[2][22] ,
         \key_mem[2][21] , \key_mem[2][20] , \key_mem[2][19] ,
         \key_mem[2][18] , \key_mem[2][17] , \key_mem[2][16] ,
         \key_mem[2][15] , \key_mem[2][14] , \key_mem[2][13] ,
         \key_mem[2][12] , \key_mem[2][11] , \key_mem[2][10] , \key_mem[2][9] ,
         \key_mem[2][8] , \key_mem[2][7] , \key_mem[2][6] , \key_mem[2][5] ,
         \key_mem[2][4] , \key_mem[2][3] , \key_mem[2][2] , \key_mem[2][1] ,
         \key_mem[2][0] , \key_mem[3][127] , \key_mem[3][126] ,
         \key_mem[3][125] , \key_mem[3][124] , \key_mem[3][123] ,
         \key_mem[3][122] , \key_mem[3][121] , \key_mem[3][120] ,
         \key_mem[3][119] , \key_mem[3][118] , \key_mem[3][117] ,
         \key_mem[3][116] , \key_mem[3][115] , \key_mem[3][114] ,
         \key_mem[3][113] , \key_mem[3][112] , \key_mem[3][111] ,
         \key_mem[3][110] , \key_mem[3][109] , \key_mem[3][108] ,
         \key_mem[3][107] , \key_mem[3][106] , \key_mem[3][105] ,
         \key_mem[3][104] , \key_mem[3][103] , \key_mem[3][102] ,
         \key_mem[3][101] , \key_mem[3][100] , \key_mem[3][99] ,
         \key_mem[3][98] , \key_mem[3][97] , \key_mem[3][96] ,
         \key_mem[3][95] , \key_mem[3][94] , \key_mem[3][93] ,
         \key_mem[3][92] , \key_mem[3][91] , \key_mem[3][90] ,
         \key_mem[3][89] , \key_mem[3][88] , \key_mem[3][87] ,
         \key_mem[3][86] , \key_mem[3][85] , \key_mem[3][84] ,
         \key_mem[3][83] , \key_mem[3][82] , \key_mem[3][81] ,
         \key_mem[3][80] , \key_mem[3][79] , \key_mem[3][78] ,
         \key_mem[3][77] , \key_mem[3][76] , \key_mem[3][75] ,
         \key_mem[3][74] , \key_mem[3][73] , \key_mem[3][72] ,
         \key_mem[3][71] , \key_mem[3][70] , \key_mem[3][69] ,
         \key_mem[3][68] , \key_mem[3][67] , \key_mem[3][66] ,
         \key_mem[3][65] , \key_mem[3][64] , \key_mem[3][63] ,
         \key_mem[3][62] , \key_mem[3][61] , \key_mem[3][60] ,
         \key_mem[3][59] , \key_mem[3][58] , \key_mem[3][57] ,
         \key_mem[3][56] , \key_mem[3][55] , \key_mem[3][54] ,
         \key_mem[3][53] , \key_mem[3][52] , \key_mem[3][51] ,
         \key_mem[3][50] , \key_mem[3][49] , \key_mem[3][48] ,
         \key_mem[3][47] , \key_mem[3][46] , \key_mem[3][45] ,
         \key_mem[3][44] , \key_mem[3][43] , \key_mem[3][42] ,
         \key_mem[3][41] , \key_mem[3][40] , \key_mem[3][39] ,
         \key_mem[3][38] , \key_mem[3][37] , \key_mem[3][36] ,
         \key_mem[3][35] , \key_mem[3][34] , \key_mem[3][33] ,
         \key_mem[3][32] , \key_mem[3][31] , \key_mem[3][30] ,
         \key_mem[3][29] , \key_mem[3][28] , \key_mem[3][27] ,
         \key_mem[3][26] , \key_mem[3][25] , \key_mem[3][24] ,
         \key_mem[3][23] , \key_mem[3][22] , \key_mem[3][21] ,
         \key_mem[3][20] , \key_mem[3][19] , \key_mem[3][18] ,
         \key_mem[3][17] , \key_mem[3][16] , \key_mem[3][15] ,
         \key_mem[3][14] , \key_mem[3][13] , \key_mem[3][12] ,
         \key_mem[3][11] , \key_mem[3][10] , \key_mem[3][9] , \key_mem[3][8] ,
         \key_mem[3][7] , \key_mem[3][6] , \key_mem[3][5] , \key_mem[3][4] ,
         \key_mem[3][3] , \key_mem[3][2] , \key_mem[3][1] , \key_mem[3][0] ,
         \key_mem[4][127] , \key_mem[4][126] , \key_mem[4][125] ,
         \key_mem[4][124] , \key_mem[4][123] , \key_mem[4][122] ,
         \key_mem[4][121] , \key_mem[4][120] , \key_mem[4][119] ,
         \key_mem[4][118] , \key_mem[4][117] , \key_mem[4][116] ,
         \key_mem[4][115] , \key_mem[4][114] , \key_mem[4][113] ,
         \key_mem[4][112] , \key_mem[4][111] , \key_mem[4][110] ,
         \key_mem[4][109] , \key_mem[4][108] , \key_mem[4][107] ,
         \key_mem[4][106] , \key_mem[4][105] , \key_mem[4][104] ,
         \key_mem[4][103] , \key_mem[4][102] , \key_mem[4][101] ,
         \key_mem[4][100] , \key_mem[4][99] , \key_mem[4][98] ,
         \key_mem[4][97] , \key_mem[4][96] , \key_mem[4][95] ,
         \key_mem[4][94] , \key_mem[4][93] , \key_mem[4][92] ,
         \key_mem[4][91] , \key_mem[4][90] , \key_mem[4][89] ,
         \key_mem[4][88] , \key_mem[4][87] , \key_mem[4][86] ,
         \key_mem[4][85] , \key_mem[4][84] , \key_mem[4][83] ,
         \key_mem[4][82] , \key_mem[4][81] , \key_mem[4][80] ,
         \key_mem[4][79] , \key_mem[4][78] , \key_mem[4][77] ,
         \key_mem[4][76] , \key_mem[4][75] , \key_mem[4][74] ,
         \key_mem[4][73] , \key_mem[4][72] , \key_mem[4][71] ,
         \key_mem[4][70] , \key_mem[4][69] , \key_mem[4][68] ,
         \key_mem[4][67] , \key_mem[4][66] , \key_mem[4][65] ,
         \key_mem[4][64] , \key_mem[4][63] , \key_mem[4][62] ,
         \key_mem[4][61] , \key_mem[4][60] , \key_mem[4][59] ,
         \key_mem[4][58] , \key_mem[4][57] , \key_mem[4][56] ,
         \key_mem[4][55] , \key_mem[4][54] , \key_mem[4][53] ,
         \key_mem[4][52] , \key_mem[4][51] , \key_mem[4][50] ,
         \key_mem[4][49] , \key_mem[4][48] , \key_mem[4][47] ,
         \key_mem[4][46] , \key_mem[4][45] , \key_mem[4][44] ,
         \key_mem[4][43] , \key_mem[4][42] , \key_mem[4][41] ,
         \key_mem[4][40] , \key_mem[4][39] , \key_mem[4][38] ,
         \key_mem[4][37] , \key_mem[4][36] , \key_mem[4][35] ,
         \key_mem[4][34] , \key_mem[4][33] , \key_mem[4][32] ,
         \key_mem[4][31] , \key_mem[4][30] , \key_mem[4][29] ,
         \key_mem[4][28] , \key_mem[4][27] , \key_mem[4][26] ,
         \key_mem[4][25] , \key_mem[4][24] , \key_mem[4][23] ,
         \key_mem[4][22] , \key_mem[4][21] , \key_mem[4][20] ,
         \key_mem[4][19] , \key_mem[4][18] , \key_mem[4][17] ,
         \key_mem[4][16] , \key_mem[4][15] , \key_mem[4][14] ,
         \key_mem[4][13] , \key_mem[4][12] , \key_mem[4][11] ,
         \key_mem[4][10] , \key_mem[4][9] , \key_mem[4][8] , \key_mem[4][7] ,
         \key_mem[4][6] , \key_mem[4][5] , \key_mem[4][4] , \key_mem[4][3] ,
         \key_mem[4][2] , \key_mem[4][1] , \key_mem[4][0] , \key_mem[5][127] ,
         \key_mem[5][126] , \key_mem[5][125] , \key_mem[5][124] ,
         \key_mem[5][123] , \key_mem[5][122] , \key_mem[5][121] ,
         \key_mem[5][120] , \key_mem[5][119] , \key_mem[5][118] ,
         \key_mem[5][117] , \key_mem[5][116] , \key_mem[5][115] ,
         \key_mem[5][114] , \key_mem[5][113] , \key_mem[5][112] ,
         \key_mem[5][111] , \key_mem[5][110] , \key_mem[5][109] ,
         \key_mem[5][108] , \key_mem[5][107] , \key_mem[5][106] ,
         \key_mem[5][105] , \key_mem[5][104] , \key_mem[5][103] ,
         \key_mem[5][102] , \key_mem[5][101] , \key_mem[5][100] ,
         \key_mem[5][99] , \key_mem[5][98] , \key_mem[5][97] ,
         \key_mem[5][96] , \key_mem[5][95] , \key_mem[5][94] ,
         \key_mem[5][93] , \key_mem[5][92] , \key_mem[5][91] ,
         \key_mem[5][90] , \key_mem[5][89] , \key_mem[5][88] ,
         \key_mem[5][87] , \key_mem[5][86] , \key_mem[5][85] ,
         \key_mem[5][84] , \key_mem[5][83] , \key_mem[5][82] ,
         \key_mem[5][81] , \key_mem[5][80] , \key_mem[5][79] ,
         \key_mem[5][78] , \key_mem[5][77] , \key_mem[5][76] ,
         \key_mem[5][75] , \key_mem[5][74] , \key_mem[5][73] ,
         \key_mem[5][72] , \key_mem[5][71] , \key_mem[5][70] ,
         \key_mem[5][69] , \key_mem[5][68] , \key_mem[5][67] ,
         \key_mem[5][66] , \key_mem[5][65] , \key_mem[5][64] ,
         \key_mem[5][63] , \key_mem[5][62] , \key_mem[5][61] ,
         \key_mem[5][60] , \key_mem[5][59] , \key_mem[5][58] ,
         \key_mem[5][57] , \key_mem[5][56] , \key_mem[5][55] ,
         \key_mem[5][54] , \key_mem[5][53] , \key_mem[5][52] ,
         \key_mem[5][51] , \key_mem[5][50] , \key_mem[5][49] ,
         \key_mem[5][48] , \key_mem[5][47] , \key_mem[5][46] ,
         \key_mem[5][45] , \key_mem[5][44] , \key_mem[5][43] ,
         \key_mem[5][42] , \key_mem[5][41] , \key_mem[5][40] ,
         \key_mem[5][39] , \key_mem[5][38] , \key_mem[5][37] ,
         \key_mem[5][36] , \key_mem[5][35] , \key_mem[5][34] ,
         \key_mem[5][33] , \key_mem[5][32] , \key_mem[5][31] ,
         \key_mem[5][30] , \key_mem[5][29] , \key_mem[5][28] ,
         \key_mem[5][27] , \key_mem[5][26] , \key_mem[5][25] ,
         \key_mem[5][24] , \key_mem[5][23] , \key_mem[5][22] ,
         \key_mem[5][21] , \key_mem[5][20] , \key_mem[5][19] ,
         \key_mem[5][18] , \key_mem[5][17] , \key_mem[5][16] ,
         \key_mem[5][15] , \key_mem[5][14] , \key_mem[5][13] ,
         \key_mem[5][12] , \key_mem[5][11] , \key_mem[5][10] , \key_mem[5][9] ,
         \key_mem[5][8] , \key_mem[5][7] , \key_mem[5][6] , \key_mem[5][5] ,
         \key_mem[5][4] , \key_mem[5][3] , \key_mem[5][2] , \key_mem[5][1] ,
         \key_mem[5][0] , \key_mem[6][127] , \key_mem[6][126] ,
         \key_mem[6][125] , \key_mem[6][124] , \key_mem[6][123] ,
         \key_mem[6][122] , \key_mem[6][121] , \key_mem[6][120] ,
         \key_mem[6][119] , \key_mem[6][118] , \key_mem[6][117] ,
         \key_mem[6][116] , \key_mem[6][115] , \key_mem[6][114] ,
         \key_mem[6][113] , \key_mem[6][112] , \key_mem[6][111] ,
         \key_mem[6][110] , \key_mem[6][109] , \key_mem[6][108] ,
         \key_mem[6][107] , \key_mem[6][106] , \key_mem[6][105] ,
         \key_mem[6][104] , \key_mem[6][103] , \key_mem[6][102] ,
         \key_mem[6][101] , \key_mem[6][100] , \key_mem[6][99] ,
         \key_mem[6][98] , \key_mem[6][97] , \key_mem[6][96] ,
         \key_mem[6][95] , \key_mem[6][94] , \key_mem[6][93] ,
         \key_mem[6][92] , \key_mem[6][91] , \key_mem[6][90] ,
         \key_mem[6][89] , \key_mem[6][88] , \key_mem[6][87] ,
         \key_mem[6][86] , \key_mem[6][85] , \key_mem[6][84] ,
         \key_mem[6][83] , \key_mem[6][82] , \key_mem[6][81] ,
         \key_mem[6][80] , \key_mem[6][79] , \key_mem[6][78] ,
         \key_mem[6][77] , \key_mem[6][76] , \key_mem[6][75] ,
         \key_mem[6][74] , \key_mem[6][73] , \key_mem[6][72] ,
         \key_mem[6][71] , \key_mem[6][70] , \key_mem[6][69] ,
         \key_mem[6][68] , \key_mem[6][67] , \key_mem[6][66] ,
         \key_mem[6][65] , \key_mem[6][64] , \key_mem[6][63] ,
         \key_mem[6][62] , \key_mem[6][61] , \key_mem[6][60] ,
         \key_mem[6][59] , \key_mem[6][58] , \key_mem[6][57] ,
         \key_mem[6][56] , \key_mem[6][55] , \key_mem[6][54] ,
         \key_mem[6][53] , \key_mem[6][52] , \key_mem[6][51] ,
         \key_mem[6][50] , \key_mem[6][49] , \key_mem[6][48] ,
         \key_mem[6][47] , \key_mem[6][46] , \key_mem[6][45] ,
         \key_mem[6][44] , \key_mem[6][43] , \key_mem[6][42] ,
         \key_mem[6][41] , \key_mem[6][40] , \key_mem[6][39] ,
         \key_mem[6][38] , \key_mem[6][37] , \key_mem[6][36] ,
         \key_mem[6][35] , \key_mem[6][34] , \key_mem[6][33] ,
         \key_mem[6][32] , \key_mem[6][31] , \key_mem[6][30] ,
         \key_mem[6][29] , \key_mem[6][28] , \key_mem[6][27] ,
         \key_mem[6][26] , \key_mem[6][25] , \key_mem[6][24] ,
         \key_mem[6][23] , \key_mem[6][22] , \key_mem[6][21] ,
         \key_mem[6][20] , \key_mem[6][19] , \key_mem[6][18] ,
         \key_mem[6][17] , \key_mem[6][16] , \key_mem[6][15] ,
         \key_mem[6][14] , \key_mem[6][13] , \key_mem[6][12] ,
         \key_mem[6][11] , \key_mem[6][10] , \key_mem[6][9] , \key_mem[6][8] ,
         \key_mem[6][7] , \key_mem[6][6] , \key_mem[6][5] , \key_mem[6][4] ,
         \key_mem[6][3] , \key_mem[6][2] , \key_mem[6][1] , \key_mem[6][0] ,
         \key_mem[7][127] , \key_mem[7][126] , \key_mem[7][125] ,
         \key_mem[7][124] , \key_mem[7][123] , \key_mem[7][122] ,
         \key_mem[7][121] , \key_mem[7][120] , \key_mem[7][119] ,
         \key_mem[7][118] , \key_mem[7][117] , \key_mem[7][116] ,
         \key_mem[7][115] , \key_mem[7][114] , \key_mem[7][113] ,
         \key_mem[7][112] , \key_mem[7][111] , \key_mem[7][110] ,
         \key_mem[7][109] , \key_mem[7][108] , \key_mem[7][107] ,
         \key_mem[7][106] , \key_mem[7][105] , \key_mem[7][104] ,
         \key_mem[7][103] , \key_mem[7][102] , \key_mem[7][101] ,
         \key_mem[7][100] , \key_mem[7][99] , \key_mem[7][98] ,
         \key_mem[7][97] , \key_mem[7][96] , \key_mem[7][95] ,
         \key_mem[7][94] , \key_mem[7][93] , \key_mem[7][92] ,
         \key_mem[7][91] , \key_mem[7][90] , \key_mem[7][89] ,
         \key_mem[7][88] , \key_mem[7][87] , \key_mem[7][86] ,
         \key_mem[7][85] , \key_mem[7][84] , \key_mem[7][83] ,
         \key_mem[7][82] , \key_mem[7][81] , \key_mem[7][80] ,
         \key_mem[7][79] , \key_mem[7][78] , \key_mem[7][77] ,
         \key_mem[7][76] , \key_mem[7][75] , \key_mem[7][74] ,
         \key_mem[7][73] , \key_mem[7][72] , \key_mem[7][71] ,
         \key_mem[7][70] , \key_mem[7][69] , \key_mem[7][68] ,
         \key_mem[7][67] , \key_mem[7][66] , \key_mem[7][65] ,
         \key_mem[7][64] , \key_mem[7][63] , \key_mem[7][62] ,
         \key_mem[7][61] , \key_mem[7][60] , \key_mem[7][59] ,
         \key_mem[7][58] , \key_mem[7][57] , \key_mem[7][56] ,
         \key_mem[7][55] , \key_mem[7][54] , \key_mem[7][53] ,
         \key_mem[7][52] , \key_mem[7][51] , \key_mem[7][50] ,
         \key_mem[7][49] , \key_mem[7][48] , \key_mem[7][47] ,
         \key_mem[7][46] , \key_mem[7][45] , \key_mem[7][44] ,
         \key_mem[7][43] , \key_mem[7][42] , \key_mem[7][41] ,
         \key_mem[7][40] , \key_mem[7][39] , \key_mem[7][38] ,
         \key_mem[7][37] , \key_mem[7][36] , \key_mem[7][35] ,
         \key_mem[7][34] , \key_mem[7][33] , \key_mem[7][32] ,
         \key_mem[7][31] , \key_mem[7][30] , \key_mem[7][29] ,
         \key_mem[7][28] , \key_mem[7][27] , \key_mem[7][26] ,
         \key_mem[7][25] , \key_mem[7][24] , \key_mem[7][23] ,
         \key_mem[7][22] , \key_mem[7][21] , \key_mem[7][20] ,
         \key_mem[7][19] , \key_mem[7][18] , \key_mem[7][17] ,
         \key_mem[7][16] , \key_mem[7][15] , \key_mem[7][14] ,
         \key_mem[7][13] , \key_mem[7][12] , \key_mem[7][11] ,
         \key_mem[7][10] , \key_mem[7][9] , \key_mem[7][8] , \key_mem[7][7] ,
         \key_mem[7][6] , \key_mem[7][5] , \key_mem[7][4] , \key_mem[7][3] ,
         \key_mem[7][2] , \key_mem[7][1] , \key_mem[7][0] , \key_mem[8][127] ,
         \key_mem[8][126] , \key_mem[8][125] , \key_mem[8][124] ,
         \key_mem[8][123] , \key_mem[8][122] , \key_mem[8][121] ,
         \key_mem[8][120] , \key_mem[8][119] , \key_mem[8][118] ,
         \key_mem[8][117] , \key_mem[8][116] , \key_mem[8][115] ,
         \key_mem[8][114] , \key_mem[8][113] , \key_mem[8][112] ,
         \key_mem[8][111] , \key_mem[8][110] , \key_mem[8][109] ,
         \key_mem[8][108] , \key_mem[8][107] , \key_mem[8][106] ,
         \key_mem[8][105] , \key_mem[8][104] , \key_mem[8][103] ,
         \key_mem[8][102] , \key_mem[8][101] , \key_mem[8][100] ,
         \key_mem[8][99] , \key_mem[8][98] , \key_mem[8][97] ,
         \key_mem[8][96] , \key_mem[8][95] , \key_mem[8][94] ,
         \key_mem[8][93] , \key_mem[8][92] , \key_mem[8][91] ,
         \key_mem[8][90] , \key_mem[8][89] , \key_mem[8][88] ,
         \key_mem[8][87] , \key_mem[8][86] , \key_mem[8][85] ,
         \key_mem[8][84] , \key_mem[8][83] , \key_mem[8][82] ,
         \key_mem[8][81] , \key_mem[8][80] , \key_mem[8][79] ,
         \key_mem[8][78] , \key_mem[8][77] , \key_mem[8][76] ,
         \key_mem[8][75] , \key_mem[8][74] , \key_mem[8][73] ,
         \key_mem[8][72] , \key_mem[8][71] , \key_mem[8][70] ,
         \key_mem[8][69] , \key_mem[8][68] , \key_mem[8][67] ,
         \key_mem[8][66] , \key_mem[8][65] , \key_mem[8][64] ,
         \key_mem[8][63] , \key_mem[8][62] , \key_mem[8][61] ,
         \key_mem[8][60] , \key_mem[8][59] , \key_mem[8][58] ,
         \key_mem[8][57] , \key_mem[8][56] , \key_mem[8][55] ,
         \key_mem[8][54] , \key_mem[8][53] , \key_mem[8][52] ,
         \key_mem[8][51] , \key_mem[8][50] , \key_mem[8][49] ,
         \key_mem[8][48] , \key_mem[8][47] , \key_mem[8][46] ,
         \key_mem[8][45] , \key_mem[8][44] , \key_mem[8][43] ,
         \key_mem[8][42] , \key_mem[8][41] , \key_mem[8][40] ,
         \key_mem[8][39] , \key_mem[8][38] , \key_mem[8][37] ,
         \key_mem[8][36] , \key_mem[8][35] , \key_mem[8][34] ,
         \key_mem[8][33] , \key_mem[8][32] , \key_mem[8][31] ,
         \key_mem[8][30] , \key_mem[8][29] , \key_mem[8][28] ,
         \key_mem[8][27] , \key_mem[8][26] , \key_mem[8][25] ,
         \key_mem[8][24] , \key_mem[8][23] , \key_mem[8][22] ,
         \key_mem[8][21] , \key_mem[8][20] , \key_mem[8][19] ,
         \key_mem[8][18] , \key_mem[8][17] , \key_mem[8][16] ,
         \key_mem[8][15] , \key_mem[8][14] , \key_mem[8][13] ,
         \key_mem[8][12] , \key_mem[8][11] , \key_mem[8][10] , \key_mem[8][9] ,
         \key_mem[8][8] , \key_mem[8][7] , \key_mem[8][6] , \key_mem[8][5] ,
         \key_mem[8][4] , \key_mem[8][3] , \key_mem[8][2] , \key_mem[8][1] ,
         \key_mem[8][0] , \key_mem[9][127] , \key_mem[9][126] ,
         \key_mem[9][125] , \key_mem[9][124] , \key_mem[9][123] ,
         \key_mem[9][122] , \key_mem[9][121] , \key_mem[9][120] ,
         \key_mem[9][119] , \key_mem[9][118] , \key_mem[9][117] ,
         \key_mem[9][116] , \key_mem[9][115] , \key_mem[9][114] ,
         \key_mem[9][113] , \key_mem[9][112] , \key_mem[9][111] ,
         \key_mem[9][110] , \key_mem[9][109] , \key_mem[9][108] ,
         \key_mem[9][107] , \key_mem[9][106] , \key_mem[9][105] ,
         \key_mem[9][104] , \key_mem[9][103] , \key_mem[9][102] ,
         \key_mem[9][101] , \key_mem[9][100] , \key_mem[9][99] ,
         \key_mem[9][98] , \key_mem[9][97] , \key_mem[9][96] ,
         \key_mem[9][95] , \key_mem[9][94] , \key_mem[9][93] ,
         \key_mem[9][92] , \key_mem[9][91] , \key_mem[9][90] ,
         \key_mem[9][89] , \key_mem[9][88] , \key_mem[9][87] ,
         \key_mem[9][86] , \key_mem[9][85] , \key_mem[9][84] ,
         \key_mem[9][83] , \key_mem[9][82] , \key_mem[9][81] ,
         \key_mem[9][80] , \key_mem[9][79] , \key_mem[9][78] ,
         \key_mem[9][77] , \key_mem[9][76] , \key_mem[9][75] ,
         \key_mem[9][74] , \key_mem[9][73] , \key_mem[9][72] ,
         \key_mem[9][71] , \key_mem[9][70] , \key_mem[9][69] ,
         \key_mem[9][68] , \key_mem[9][67] , \key_mem[9][66] ,
         \key_mem[9][65] , \key_mem[9][64] , \key_mem[9][63] ,
         \key_mem[9][62] , \key_mem[9][61] , \key_mem[9][60] ,
         \key_mem[9][59] , \key_mem[9][58] , \key_mem[9][57] ,
         \key_mem[9][56] , \key_mem[9][55] , \key_mem[9][54] ,
         \key_mem[9][53] , \key_mem[9][52] , \key_mem[9][51] ,
         \key_mem[9][50] , \key_mem[9][49] , \key_mem[9][48] ,
         \key_mem[9][47] , \key_mem[9][46] , \key_mem[9][45] ,
         \key_mem[9][44] , \key_mem[9][43] , \key_mem[9][42] ,
         \key_mem[9][41] , \key_mem[9][40] , \key_mem[9][39] ,
         \key_mem[9][38] , \key_mem[9][37] , \key_mem[9][36] ,
         \key_mem[9][35] , \key_mem[9][34] , \key_mem[9][33] ,
         \key_mem[9][32] , \key_mem[9][31] , \key_mem[9][30] ,
         \key_mem[9][29] , \key_mem[9][28] , \key_mem[9][27] ,
         \key_mem[9][26] , \key_mem[9][25] , \key_mem[9][24] ,
         \key_mem[9][23] , \key_mem[9][22] , \key_mem[9][21] ,
         \key_mem[9][20] , \key_mem[9][19] , \key_mem[9][18] ,
         \key_mem[9][17] , \key_mem[9][16] , \key_mem[9][15] ,
         \key_mem[9][14] , \key_mem[9][13] , \key_mem[9][12] ,
         \key_mem[9][11] , \key_mem[9][10] , \key_mem[9][9] , \key_mem[9][8] ,
         \key_mem[9][7] , \key_mem[9][6] , \key_mem[9][5] , \key_mem[9][4] ,
         \key_mem[9][3] , \key_mem[9][2] , \key_mem[9][1] , \key_mem[9][0] ,
         \key_mem[10][127] , \key_mem[10][126] , \key_mem[10][125] ,
         \key_mem[10][124] , \key_mem[10][123] , \key_mem[10][122] ,
         \key_mem[10][121] , \key_mem[10][120] , \key_mem[10][119] ,
         \key_mem[10][118] , \key_mem[10][117] , \key_mem[10][116] ,
         \key_mem[10][115] , \key_mem[10][114] , \key_mem[10][113] ,
         \key_mem[10][112] , \key_mem[10][111] , \key_mem[10][110] ,
         \key_mem[10][109] , \key_mem[10][108] , \key_mem[10][107] ,
         \key_mem[10][106] , \key_mem[10][105] , \key_mem[10][104] ,
         \key_mem[10][103] , \key_mem[10][102] , \key_mem[10][101] ,
         \key_mem[10][100] , \key_mem[10][99] , \key_mem[10][98] ,
         \key_mem[10][97] , \key_mem[10][96] , \key_mem[10][95] ,
         \key_mem[10][94] , \key_mem[10][93] , \key_mem[10][92] ,
         \key_mem[10][91] , \key_mem[10][90] , \key_mem[10][89] ,
         \key_mem[10][88] , \key_mem[10][87] , \key_mem[10][86] ,
         \key_mem[10][85] , \key_mem[10][84] , \key_mem[10][83] ,
         \key_mem[10][82] , \key_mem[10][81] , \key_mem[10][80] ,
         \key_mem[10][79] , \key_mem[10][78] , \key_mem[10][77] ,
         \key_mem[10][76] , \key_mem[10][75] , \key_mem[10][74] ,
         \key_mem[10][73] , \key_mem[10][72] , \key_mem[10][71] ,
         \key_mem[10][70] , \key_mem[10][69] , \key_mem[10][68] ,
         \key_mem[10][67] , \key_mem[10][66] , \key_mem[10][65] ,
         \key_mem[10][64] , \key_mem[10][63] , \key_mem[10][62] ,
         \key_mem[10][61] , \key_mem[10][60] , \key_mem[10][59] ,
         \key_mem[10][58] , \key_mem[10][57] , \key_mem[10][56] ,
         \key_mem[10][55] , \key_mem[10][54] , \key_mem[10][53] ,
         \key_mem[10][52] , \key_mem[10][51] , \key_mem[10][50] ,
         \key_mem[10][49] , \key_mem[10][48] , \key_mem[10][47] ,
         \key_mem[10][46] , \key_mem[10][45] , \key_mem[10][44] ,
         \key_mem[10][43] , \key_mem[10][42] , \key_mem[10][41] ,
         \key_mem[10][40] , \key_mem[10][39] , \key_mem[10][38] ,
         \key_mem[10][37] , \key_mem[10][36] , \key_mem[10][35] ,
         \key_mem[10][34] , \key_mem[10][33] , \key_mem[10][32] ,
         \key_mem[10][31] , \key_mem[10][30] , \key_mem[10][29] ,
         \key_mem[10][28] , \key_mem[10][27] , \key_mem[10][26] ,
         \key_mem[10][25] , \key_mem[10][24] , \key_mem[10][23] ,
         \key_mem[10][22] , \key_mem[10][21] , \key_mem[10][20] ,
         \key_mem[10][19] , \key_mem[10][18] , \key_mem[10][17] ,
         \key_mem[10][16] , \key_mem[10][15] , \key_mem[10][14] ,
         \key_mem[10][13] , \key_mem[10][12] , \key_mem[10][11] ,
         \key_mem[10][10] , \key_mem[10][9] , \key_mem[10][8] ,
         \key_mem[10][7] , \key_mem[10][6] , \key_mem[10][5] ,
         \key_mem[10][4] , \key_mem[10][3] , \key_mem[10][2] ,
         \key_mem[10][1] , \key_mem[10][0] , \key_mem[11][127] ,
         \key_mem[11][126] , \key_mem[11][125] , \key_mem[11][124] ,
         \key_mem[11][123] , \key_mem[11][122] , \key_mem[11][121] ,
         \key_mem[11][120] , \key_mem[11][119] , \key_mem[11][118] ,
         \key_mem[11][117] , \key_mem[11][116] , \key_mem[11][115] ,
         \key_mem[11][114] , \key_mem[11][113] , \key_mem[11][112] ,
         \key_mem[11][111] , \key_mem[11][110] , \key_mem[11][109] ,
         \key_mem[11][108] , \key_mem[11][107] , \key_mem[11][106] ,
         \key_mem[11][105] , \key_mem[11][104] , \key_mem[11][103] ,
         \key_mem[11][102] , \key_mem[11][101] , \key_mem[11][100] ,
         \key_mem[11][99] , \key_mem[11][98] , \key_mem[11][97] ,
         \key_mem[11][96] , \key_mem[11][95] , \key_mem[11][94] ,
         \key_mem[11][93] , \key_mem[11][92] , \key_mem[11][91] ,
         \key_mem[11][90] , \key_mem[11][89] , \key_mem[11][88] ,
         \key_mem[11][87] , \key_mem[11][86] , \key_mem[11][85] ,
         \key_mem[11][84] , \key_mem[11][83] , \key_mem[11][82] ,
         \key_mem[11][81] , \key_mem[11][80] , \key_mem[11][79] ,
         \key_mem[11][78] , \key_mem[11][77] , \key_mem[11][76] ,
         \key_mem[11][75] , \key_mem[11][74] , \key_mem[11][73] ,
         \key_mem[11][72] , \key_mem[11][71] , \key_mem[11][70] ,
         \key_mem[11][69] , \key_mem[11][68] , \key_mem[11][67] ,
         \key_mem[11][66] , \key_mem[11][65] , \key_mem[11][64] ,
         \key_mem[11][63] , \key_mem[11][62] , \key_mem[11][61] ,
         \key_mem[11][60] , \key_mem[11][59] , \key_mem[11][58] ,
         \key_mem[11][57] , \key_mem[11][56] , \key_mem[11][55] ,
         \key_mem[11][54] , \key_mem[11][53] , \key_mem[11][52] ,
         \key_mem[11][51] , \key_mem[11][50] , \key_mem[11][49] ,
         \key_mem[11][48] , \key_mem[11][47] , \key_mem[11][46] ,
         \key_mem[11][45] , \key_mem[11][44] , \key_mem[11][43] ,
         \key_mem[11][42] , \key_mem[11][41] , \key_mem[11][40] ,
         \key_mem[11][39] , \key_mem[11][38] , \key_mem[11][37] ,
         \key_mem[11][36] , \key_mem[11][35] , \key_mem[11][34] ,
         \key_mem[11][33] , \key_mem[11][32] , \key_mem[11][31] ,
         \key_mem[11][30] , \key_mem[11][29] , \key_mem[11][28] ,
         \key_mem[11][27] , \key_mem[11][26] , \key_mem[11][25] ,
         \key_mem[11][24] , \key_mem[11][23] , \key_mem[11][22] ,
         \key_mem[11][21] , \key_mem[11][20] , \key_mem[11][19] ,
         \key_mem[11][18] , \key_mem[11][17] , \key_mem[11][16] ,
         \key_mem[11][15] , \key_mem[11][14] , \key_mem[11][13] ,
         \key_mem[11][12] , \key_mem[11][11] , \key_mem[11][10] ,
         \key_mem[11][9] , \key_mem[11][8] , \key_mem[11][7] ,
         \key_mem[11][6] , \key_mem[11][5] , \key_mem[11][4] ,
         \key_mem[11][3] , \key_mem[11][2] , \key_mem[11][1] ,
         \key_mem[11][0] , \key_mem[12][127] , \key_mem[12][126] ,
         \key_mem[12][125] , \key_mem[12][124] , \key_mem[12][123] ,
         \key_mem[12][122] , \key_mem[12][121] , \key_mem[12][120] ,
         \key_mem[12][119] , \key_mem[12][118] , \key_mem[12][117] ,
         \key_mem[12][116] , \key_mem[12][115] , \key_mem[12][114] ,
         \key_mem[12][113] , \key_mem[12][112] , \key_mem[12][111] ,
         \key_mem[12][110] , \key_mem[12][109] , \key_mem[12][108] ,
         \key_mem[12][107] , \key_mem[12][106] , \key_mem[12][105] ,
         \key_mem[12][104] , \key_mem[12][103] , \key_mem[12][102] ,
         \key_mem[12][101] , \key_mem[12][100] , \key_mem[12][99] ,
         \key_mem[12][98] , \key_mem[12][97] , \key_mem[12][96] ,
         \key_mem[12][95] , \key_mem[12][94] , \key_mem[12][93] ,
         \key_mem[12][92] , \key_mem[12][91] , \key_mem[12][90] ,
         \key_mem[12][89] , \key_mem[12][88] , \key_mem[12][87] ,
         \key_mem[12][86] , \key_mem[12][85] , \key_mem[12][84] ,
         \key_mem[12][83] , \key_mem[12][82] , \key_mem[12][81] ,
         \key_mem[12][80] , \key_mem[12][79] , \key_mem[12][78] ,
         \key_mem[12][77] , \key_mem[12][76] , \key_mem[12][75] ,
         \key_mem[12][74] , \key_mem[12][73] , \key_mem[12][72] ,
         \key_mem[12][71] , \key_mem[12][70] , \key_mem[12][69] ,
         \key_mem[12][68] , \key_mem[12][67] , \key_mem[12][66] ,
         \key_mem[12][65] , \key_mem[12][64] , \key_mem[12][63] ,
         \key_mem[12][62] , \key_mem[12][61] , \key_mem[12][60] ,
         \key_mem[12][59] , \key_mem[12][58] , \key_mem[12][57] ,
         \key_mem[12][56] , \key_mem[12][55] , \key_mem[12][54] ,
         \key_mem[12][53] , \key_mem[12][52] , \key_mem[12][51] ,
         \key_mem[12][50] , \key_mem[12][49] , \key_mem[12][48] ,
         \key_mem[12][47] , \key_mem[12][46] , \key_mem[12][45] ,
         \key_mem[12][44] , \key_mem[12][43] , \key_mem[12][42] ,
         \key_mem[12][41] , \key_mem[12][40] , \key_mem[12][39] ,
         \key_mem[12][38] , \key_mem[12][37] , \key_mem[12][36] ,
         \key_mem[12][35] , \key_mem[12][34] , \key_mem[12][33] ,
         \key_mem[12][32] , \key_mem[12][31] , \key_mem[12][30] ,
         \key_mem[12][29] , \key_mem[12][28] , \key_mem[12][27] ,
         \key_mem[12][26] , \key_mem[12][25] , \key_mem[12][24] ,
         \key_mem[12][23] , \key_mem[12][22] , \key_mem[12][21] ,
         \key_mem[12][20] , \key_mem[12][19] , \key_mem[12][18] ,
         \key_mem[12][17] , \key_mem[12][16] , \key_mem[12][15] ,
         \key_mem[12][14] , \key_mem[12][13] , \key_mem[12][12] ,
         \key_mem[12][11] , \key_mem[12][10] , \key_mem[12][9] ,
         \key_mem[12][8] , \key_mem[12][7] , \key_mem[12][6] ,
         \key_mem[12][5] , \key_mem[12][4] , \key_mem[12][3] ,
         \key_mem[12][2] , \key_mem[12][1] , \key_mem[12][0] ,
         \key_mem[13][127] , \key_mem[13][126] , \key_mem[13][125] ,
         \key_mem[13][124] , \key_mem[13][123] , \key_mem[13][122] ,
         \key_mem[13][121] , \key_mem[13][120] , \key_mem[13][119] ,
         \key_mem[13][118] , \key_mem[13][117] , \key_mem[13][116] ,
         \key_mem[13][115] , \key_mem[13][114] , \key_mem[13][113] ,
         \key_mem[13][112] , \key_mem[13][111] , \key_mem[13][110] ,
         \key_mem[13][109] , \key_mem[13][108] , \key_mem[13][107] ,
         \key_mem[13][106] , \key_mem[13][105] , \key_mem[13][104] ,
         \key_mem[13][103] , \key_mem[13][102] , \key_mem[13][101] ,
         \key_mem[13][100] , \key_mem[13][99] , \key_mem[13][98] ,
         \key_mem[13][97] , \key_mem[13][96] , \key_mem[13][95] ,
         \key_mem[13][94] , \key_mem[13][93] , \key_mem[13][92] ,
         \key_mem[13][91] , \key_mem[13][90] , \key_mem[13][89] ,
         \key_mem[13][88] , \key_mem[13][87] , \key_mem[13][86] ,
         \key_mem[13][85] , \key_mem[13][84] , \key_mem[13][83] ,
         \key_mem[13][82] , \key_mem[13][81] , \key_mem[13][80] ,
         \key_mem[13][79] , \key_mem[13][78] , \key_mem[13][77] ,
         \key_mem[13][76] , \key_mem[13][75] , \key_mem[13][74] ,
         \key_mem[13][73] , \key_mem[13][72] , \key_mem[13][71] ,
         \key_mem[13][70] , \key_mem[13][69] , \key_mem[13][68] ,
         \key_mem[13][67] , \key_mem[13][66] , \key_mem[13][65] ,
         \key_mem[13][64] , \key_mem[13][63] , \key_mem[13][62] ,
         \key_mem[13][61] , \key_mem[13][60] , \key_mem[13][59] ,
         \key_mem[13][58] , \key_mem[13][57] , \key_mem[13][56] ,
         \key_mem[13][55] , \key_mem[13][54] , \key_mem[13][53] ,
         \key_mem[13][52] , \key_mem[13][51] , \key_mem[13][50] ,
         \key_mem[13][49] , \key_mem[13][48] , \key_mem[13][47] ,
         \key_mem[13][46] , \key_mem[13][45] , \key_mem[13][44] ,
         \key_mem[13][43] , \key_mem[13][42] , \key_mem[13][41] ,
         \key_mem[13][40] , \key_mem[13][39] , \key_mem[13][38] ,
         \key_mem[13][37] , \key_mem[13][36] , \key_mem[13][35] ,
         \key_mem[13][34] , \key_mem[13][33] , \key_mem[13][32] ,
         \key_mem[13][31] , \key_mem[13][30] , \key_mem[13][29] ,
         \key_mem[13][28] , \key_mem[13][27] , \key_mem[13][26] ,
         \key_mem[13][25] , \key_mem[13][24] , \key_mem[13][23] ,
         \key_mem[13][22] , \key_mem[13][21] , \key_mem[13][20] ,
         \key_mem[13][19] , \key_mem[13][18] , \key_mem[13][17] ,
         \key_mem[13][16] , \key_mem[13][15] , \key_mem[13][14] ,
         \key_mem[13][13] , \key_mem[13][12] , \key_mem[13][11] ,
         \key_mem[13][10] , \key_mem[13][9] , \key_mem[13][8] ,
         \key_mem[13][7] , \key_mem[13][6] , \key_mem[13][5] ,
         \key_mem[13][4] , \key_mem[13][3] , \key_mem[13][2] ,
         \key_mem[13][1] , \key_mem[13][0] , \key_mem[14][127] ,
         \key_mem[14][126] , \key_mem[14][125] , \key_mem[14][124] ,
         \key_mem[14][123] , \key_mem[14][122] , \key_mem[14][121] ,
         \key_mem[14][120] , \key_mem[14][119] , \key_mem[14][118] ,
         \key_mem[14][117] , \key_mem[14][116] , \key_mem[14][115] ,
         \key_mem[14][114] , \key_mem[14][113] , \key_mem[14][112] ,
         \key_mem[14][111] , \key_mem[14][110] , \key_mem[14][109] ,
         \key_mem[14][108] , \key_mem[14][107] , \key_mem[14][106] ,
         \key_mem[14][105] , \key_mem[14][104] , \key_mem[14][103] ,
         \key_mem[14][102] , \key_mem[14][101] , \key_mem[14][100] ,
         \key_mem[14][99] , \key_mem[14][98] , \key_mem[14][97] ,
         \key_mem[14][96] , \key_mem[14][95] , \key_mem[14][94] ,
         \key_mem[14][93] , \key_mem[14][92] , \key_mem[14][91] ,
         \key_mem[14][90] , \key_mem[14][89] , \key_mem[14][88] ,
         \key_mem[14][87] , \key_mem[14][86] , \key_mem[14][85] ,
         \key_mem[14][84] , \key_mem[14][83] , \key_mem[14][82] ,
         \key_mem[14][81] , \key_mem[14][80] , \key_mem[14][79] ,
         \key_mem[14][78] , \key_mem[14][77] , \key_mem[14][76] ,
         \key_mem[14][75] , \key_mem[14][74] , \key_mem[14][73] ,
         \key_mem[14][72] , \key_mem[14][71] , \key_mem[14][70] ,
         \key_mem[14][69] , \key_mem[14][68] , \key_mem[14][67] ,
         \key_mem[14][66] , \key_mem[14][65] , \key_mem[14][64] ,
         \key_mem[14][63] , \key_mem[14][62] , \key_mem[14][61] ,
         \key_mem[14][60] , \key_mem[14][59] , \key_mem[14][58] ,
         \key_mem[14][57] , \key_mem[14][56] , \key_mem[14][55] ,
         \key_mem[14][54] , \key_mem[14][53] , \key_mem[14][52] ,
         \key_mem[14][51] , \key_mem[14][50] , \key_mem[14][49] ,
         \key_mem[14][48] , \key_mem[14][47] , \key_mem[14][46] ,
         \key_mem[14][45] , \key_mem[14][44] , \key_mem[14][43] ,
         \key_mem[14][42] , \key_mem[14][41] , \key_mem[14][40] ,
         \key_mem[14][39] , \key_mem[14][38] , \key_mem[14][37] ,
         \key_mem[14][36] , \key_mem[14][35] , \key_mem[14][34] ,
         \key_mem[14][33] , \key_mem[14][32] , \key_mem[14][31] ,
         \key_mem[14][30] , \key_mem[14][29] , \key_mem[14][28] ,
         \key_mem[14][27] , \key_mem[14][26] , \key_mem[14][25] ,
         \key_mem[14][24] , \key_mem[14][23] , \key_mem[14][22] ,
         \key_mem[14][21] , \key_mem[14][20] , \key_mem[14][19] ,
         \key_mem[14][18] , \key_mem[14][17] , \key_mem[14][16] ,
         \key_mem[14][15] , \key_mem[14][14] , \key_mem[14][13] ,
         \key_mem[14][12] , \key_mem[14][11] , \key_mem[14][10] ,
         \key_mem[14][9] , \key_mem[14][8] , \key_mem[14][7] ,
         \key_mem[14][6] , \key_mem[14][5] , \key_mem[14][4] ,
         \key_mem[14][3] , \key_mem[14][2] , \key_mem[14][1] ,
         \key_mem[14][0] , n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n276, n277, n278, n279, n281, n283,
         n285, n287, n289, n291, n293, n295, n298, n299, n590, n591, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n749, n750, n752, n753, n754,
         n756, n757, n758, n760, n761, n762, n764, n765, n766, n768, n769,
         n770, n772, n773, n774, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n909, n910, n913, n914, n917, n918, n921, n922, n925, n926,
         n929, n930, n933, n934, n937, n938, n941, n942, n945, n946, n949,
         n950, n953, n954, n957, n958, n961, n962, n965, n966, n969, n970,
         n973, n974, n977, n978, n981, n982, n985, n986, n989, n990, n993,
         n994, n997, n998, n1001, n1002, n1005, n1006, n1008, n1009, n1010,
         n1012, n1013, n1014, n1016, n1017, n1018, n1020, n1021, n1022, n1024,
         n1025, n1026, n1028, n1029, n1030, n1032, n1033, n1034, n1035, n1037,
         n1038, n1039, n1041, n1042, n1043, n1045, n1046, n1047, n1049, n1050,
         n1051, n1053, n1054, n1055, n1057, n1058, n1059, n1061, n1062, n1063,
         n1065, n1066, n1067, n1069, n1070, n1071, n1073, n1074, n1075, n1077,
         n1078, n1079, n1081, n1082, n1083, n1085, n1086, n1087, n1089, n1090,
         n1091, n1093, n1094, n1095, n1097, n1098, n1099, n1101, n1102, n1103,
         n1105, n1106, n1107, n1109, n1110, n1111, n1113, n1114, n1115, n1117,
         n1118, n1119, n1121, n1122, n1123, n1126, n1127, n1129, n1130, n1133,
         n1134, n1136, n1137, n1138, n1140, n1141, n1142, n1144, n1145, n1146,
         n1148, n1149, n1150, n1152, n1153, n1154, n1156, n1157, n1158, n1160,
         n1161, n1162, n1165, n1166, n1169, n1170, n1173, n1174, n1177, n1178,
         n1181, n1182, n1185, n1186, n1189, n1190, n1193, n1194, n1197, n1198,
         n1201, n1202, n1205, n1206, n1209, n1210, n1213, n1214, n1217, n1218,
         n1221, n1222, n1225, n1226, n1229, n1230, n1233, n1234, n1237, n1238,
         n1241, n1242, n1245, n1246, n1249, n1250, n1254, n1718, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n280, n282, n284, n286, n288, n290, n292, n294, n296, n297,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n592, n721, n744, n745, n746, n747, n748,
         n751, n755, n759, n763, n767, n771, n775, n875, n876, n907, n908,
         n911, n912, n915, n916, n919, n920, n923, n924, n927, n928, n931,
         n932, n935, n936, n939, n940, n943, n944, n947, n948, n951, n952,
         n955, n956, n959, n960, n963, n964, n967, n968, n971, n972, n975,
         n976, n979, n980, n983, n984, n987, n988, n991, n992, n995, n996,
         n999, n1000, n1003, n1004, n1007, n1011, n1015, n1019, n1023, n1027,
         n1031, n1036, n1040, n1044, n1048, n1052, n1056, n1060, n1064, n1068,
         n1072, n1076, n1080, n1084, n1088, n1092, n1096, n1100, n1104, n1108,
         n1112, n1116, n1120, n1124, n1125, n1128, n1131, n1132, n1135, n1139,
         n1143, n1147, n1151, n1155, n1159, n1163, n1164, n1167, n1168, n1171,
         n1172, n1175, n1176, n1179, n1180, n1183, n1184, n1187, n1188, n1191,
         n1192, n1195, n1196, n1199, n1200, n1203, n1204, n1207, n1208, n1211,
         n1212, n1215, n1216, n1219, n1220, n1223, n1224, n1227, n1228, n1231,
         n1232, n1235, n1236, n1239, n1240, n1243, n1244, n1247, n1248, n1251,
         n1252, n1253, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1719, n1720, n1728, n1736, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893;
  wire   [7:0] rcon_reg;
  wire   [2:0] key_mem_ctrl_reg;
  wire   [3:0] round_ctr_reg;
  wire   [127:0] prev_key0_reg;
  wire   [127:32] prev_key1_reg;
  assign N31 = round[0];
  assign N32 = round[1];
  assign N33 = round[2];
  assign N34 = round[3];

  DFFQX1 \prev_key0_reg_reg[105]  ( .D(n3680), .CK(clk), .Q(prev_key0_reg[105]) );
  DFFQX1 \prev_key0_reg_reg[22]  ( .D(n3762), .CK(clk), .Q(prev_key0_reg[22])
         );
  DFFQX1 \prev_key0_reg_reg[20]  ( .D(n3764), .CK(clk), .Q(prev_key0_reg[20])
         );
  DFFQX1 \prev_key0_reg_reg[17]  ( .D(n3767), .CK(clk), .Q(prev_key0_reg[17])
         );
  DFFQX1 \prev_key0_reg_reg[16]  ( .D(n3768), .CK(clk), .Q(prev_key0_reg[16])
         );
  DFFQX1 \prev_key0_reg_reg[12]  ( .D(n3772), .CK(clk), .Q(prev_key0_reg[12])
         );
  DFFQX1 \prev_key0_reg_reg[9]  ( .D(n3775), .CK(clk), .Q(prev_key0_reg[9]) );
  DFFQX1 \prev_key0_reg_reg[116]  ( .D(n3669), .CK(clk), .Q(prev_key0_reg[116]) );
  DFFQX1 \prev_key0_reg_reg[112]  ( .D(n3673), .CK(clk), .Q(prev_key0_reg[112]) );
  DFFQX1 \prev_key0_reg_reg[108]  ( .D(n3677), .CK(clk), .Q(prev_key0_reg[108]) );
  DFFQX1 \prev_key1_reg_reg[32]  ( .D(n3880), .CK(clk), .Q(prev_key1_reg[32])
         );
  DFFQX1 \prev_key1_reg_reg[44]  ( .D(n3868), .CK(clk), .Q(prev_key1_reg[44])
         );
  DFFQX1 \prev_key1_reg_reg[40]  ( .D(n3872), .CK(clk), .Q(prev_key1_reg[40])
         );
  DFFQX1 \prev_key1_reg_reg[33]  ( .D(n3879), .CK(clk), .Q(prev_key1_reg[33])
         );
  DFFQX1 \prev_key1_reg_reg[55]  ( .D(n3857), .CK(clk), .Q(prev_key1_reg[55])
         );
  DFFQX1 \prev_key1_reg_reg[54]  ( .D(n3858), .CK(clk), .Q(prev_key1_reg[54])
         );
  DFFQX1 \prev_key1_reg_reg[53]  ( .D(n3859), .CK(clk), .Q(prev_key1_reg[53])
         );
  DFFQX1 \prev_key1_reg_reg[52]  ( .D(n3860), .CK(clk), .Q(prev_key1_reg[52])
         );
  DFFQX1 \prev_key1_reg_reg[51]  ( .D(n3861), .CK(clk), .Q(prev_key1_reg[51])
         );
  DFFQX1 \prev_key1_reg_reg[50]  ( .D(n3862), .CK(clk), .Q(prev_key1_reg[50])
         );
  DFFQX1 \prev_key1_reg_reg[49]  ( .D(n3863), .CK(clk), .Q(prev_key1_reg[49])
         );
  DFFQX1 \prev_key1_reg_reg[48]  ( .D(n3864), .CK(clk), .Q(prev_key1_reg[48])
         );
  DFFQX1 \prev_key1_reg_reg[47]  ( .D(n3865), .CK(clk), .Q(prev_key1_reg[47])
         );
  DFFQX1 \prev_key1_reg_reg[46]  ( .D(n3866), .CK(clk), .Q(prev_key1_reg[46])
         );
  DFFQX1 \prev_key1_reg_reg[45]  ( .D(n3867), .CK(clk), .Q(prev_key1_reg[45])
         );
  DFFQX1 \prev_key1_reg_reg[43]  ( .D(n3869), .CK(clk), .Q(prev_key1_reg[43])
         );
  DFFQX1 \prev_key1_reg_reg[42]  ( .D(n3870), .CK(clk), .Q(prev_key1_reg[42])
         );
  DFFQX1 \prev_key1_reg_reg[41]  ( .D(n3871), .CK(clk), .Q(prev_key1_reg[41])
         );
  DFFQX1 \prev_key1_reg_reg[39]  ( .D(n3873), .CK(clk), .Q(prev_key1_reg[39])
         );
  DFFQX1 \prev_key1_reg_reg[38]  ( .D(n3874), .CK(clk), .Q(prev_key1_reg[38])
         );
  DFFQX1 \prev_key1_reg_reg[37]  ( .D(n3875), .CK(clk), .Q(prev_key1_reg[37])
         );
  DFFQX1 \prev_key1_reg_reg[36]  ( .D(n3876), .CK(clk), .Q(prev_key1_reg[36])
         );
  DFFQX1 \prev_key1_reg_reg[35]  ( .D(n3877), .CK(clk), .Q(prev_key1_reg[35])
         );
  DFFQX1 \prev_key1_reg_reg[34]  ( .D(n3878), .CK(clk), .Q(prev_key1_reg[34])
         );
  DFFQX1 \prev_key0_reg_reg[118]  ( .D(n3667), .CK(clk), .Q(prev_key0_reg[118]) );
  DFFQX1 \prev_key1_reg_reg[108]  ( .D(n3804), .CK(clk), .Q(prev_key1_reg[108]) );
  DFFQX1 \prev_key1_reg_reg[118]  ( .D(n3794), .CK(clk), .Q(prev_key1_reg[118]) );
  DFFQX1 \prev_key1_reg_reg[127]  ( .D(n3785), .CK(clk), .Q(prev_key1_reg[127]) );
  DFFQX1 \prev_key1_reg_reg[95]  ( .D(n3817), .CK(clk), .Q(prev_key1_reg[95])
         );
  DFFQX1 \prev_key1_reg_reg[63]  ( .D(n3849), .CK(clk), .Q(prev_key1_reg[63])
         );
  DFFQX1 \prev_key1_reg_reg[56]  ( .D(n3856), .CK(clk), .Q(prev_key1_reg[56])
         );
  DFFQX1 \prev_key1_reg_reg[58]  ( .D(n3854), .CK(clk), .Q(prev_key1_reg[58])
         );
  DFFQX1 \prev_key1_reg_reg[59]  ( .D(n3853), .CK(clk), .Q(prev_key1_reg[59])
         );
  DFFQX1 \prev_key1_reg_reg[62]  ( .D(n3850), .CK(clk), .Q(prev_key1_reg[62])
         );
  DFFQX1 \prev_key1_reg_reg[61]  ( .D(n3851), .CK(clk), .Q(prev_key1_reg[61])
         );
  DFFQX1 \prev_key1_reg_reg[60]  ( .D(n3852), .CK(clk), .Q(prev_key1_reg[60])
         );
  DFFQX1 \prev_key1_reg_reg[57]  ( .D(n3855), .CK(clk), .Q(prev_key1_reg[57])
         );
  DFFQX1 \prev_key0_reg_reg[54]  ( .D(n3730), .CK(clk), .Q(prev_key0_reg[54])
         );
  DFFQX1 \prev_key0_reg_reg[52]  ( .D(n3732), .CK(clk), .Q(prev_key0_reg[52])
         );
  DFFQX1 \prev_key0_reg_reg[49]  ( .D(n3735), .CK(clk), .Q(prev_key0_reg[49])
         );
  DFFQX1 \prev_key0_reg_reg[48]  ( .D(n3736), .CK(clk), .Q(prev_key0_reg[48])
         );
  DFFQX1 \prev_key0_reg_reg[44]  ( .D(n3740), .CK(clk), .Q(prev_key0_reg[44])
         );
  DFFQX1 \prev_key0_reg_reg[41]  ( .D(n3743), .CK(clk), .Q(prev_key0_reg[41])
         );
  DFFQX1 \prev_key0_reg_reg[40]  ( .D(n3744), .CK(clk), .Q(prev_key0_reg[40])
         );
  DFFQX1 \prev_key0_reg_reg[39]  ( .D(n3745), .CK(clk), .Q(prev_key0_reg[39])
         );
  DFFQX1 \prev_key0_reg_reg[38]  ( .D(n3746), .CK(clk), .Q(prev_key0_reg[38])
         );
  DFFQX1 \prev_key0_reg_reg[37]  ( .D(n3747), .CK(clk), .Q(prev_key0_reg[37])
         );
  DFFQX1 \prev_key0_reg_reg[36]  ( .D(n3748), .CK(clk), .Q(prev_key0_reg[36])
         );
  DFFQX1 \prev_key0_reg_reg[35]  ( .D(n3749), .CK(clk), .Q(prev_key0_reg[35])
         );
  DFFQX1 \prev_key0_reg_reg[34]  ( .D(n3750), .CK(clk), .Q(prev_key0_reg[34])
         );
  DFFQX1 \prev_key0_reg_reg[33]  ( .D(n3751), .CK(clk), .Q(prev_key0_reg[33])
         );
  DFFQX1 \prev_key0_reg_reg[32]  ( .D(n3752), .CK(clk), .Q(prev_key0_reg[32])
         );
  DFFQX1 \prev_key0_reg_reg[63]  ( .D(n3721), .CK(clk), .Q(prev_key0_reg[63])
         );
  DFFQX1 \prev_key1_reg_reg[78]  ( .D(n3834), .CK(clk), .Q(prev_key1_reg[78])
         );
  DFFQX1 \prev_key1_reg_reg[76]  ( .D(n3836), .CK(clk), .Q(prev_key1_reg[76])
         );
  DFFQX1 \prev_key1_reg_reg[72]  ( .D(n3840), .CK(clk), .Q(prev_key1_reg[72])
         );
  DFFQX1 \prev_key1_reg_reg[64]  ( .D(n3848), .CK(clk), .Q(prev_key1_reg[64])
         );
  DFFQX1 \prev_key1_reg_reg[68]  ( .D(n3844), .CK(clk), .Q(prev_key1_reg[68])
         );
  DFFQX1 \prev_key1_reg_reg[65]  ( .D(n3847), .CK(clk), .Q(prev_key1_reg[65])
         );
  DFFQX1 \prev_key1_reg_reg[87]  ( .D(n3825), .CK(clk), .Q(prev_key1_reg[87])
         );
  DFFQX1 \prev_key1_reg_reg[86]  ( .D(n3826), .CK(clk), .Q(prev_key1_reg[86])
         );
  DFFQX1 \prev_key1_reg_reg[85]  ( .D(n3827), .CK(clk), .Q(prev_key1_reg[85])
         );
  DFFQX1 \prev_key1_reg_reg[84]  ( .D(n3828), .CK(clk), .Q(prev_key1_reg[84])
         );
  DFFQX1 \prev_key1_reg_reg[83]  ( .D(n3829), .CK(clk), .Q(prev_key1_reg[83])
         );
  DFFQX1 \prev_key1_reg_reg[82]  ( .D(n3830), .CK(clk), .Q(prev_key1_reg[82])
         );
  DFFQX1 \prev_key1_reg_reg[81]  ( .D(n3831), .CK(clk), .Q(prev_key1_reg[81])
         );
  DFFQX1 \prev_key1_reg_reg[80]  ( .D(n3832), .CK(clk), .Q(prev_key1_reg[80])
         );
  DFFQX1 \prev_key1_reg_reg[79]  ( .D(n3833), .CK(clk), .Q(prev_key1_reg[79])
         );
  DFFQX1 \prev_key1_reg_reg[77]  ( .D(n3835), .CK(clk), .Q(prev_key1_reg[77])
         );
  DFFQX1 \prev_key1_reg_reg[75]  ( .D(n3837), .CK(clk), .Q(prev_key1_reg[75])
         );
  DFFQX1 \prev_key1_reg_reg[74]  ( .D(n3838), .CK(clk), .Q(prev_key1_reg[74])
         );
  DFFQX1 \prev_key1_reg_reg[73]  ( .D(n3839), .CK(clk), .Q(prev_key1_reg[73])
         );
  DFFQX1 \prev_key1_reg_reg[71]  ( .D(n3841), .CK(clk), .Q(prev_key1_reg[71])
         );
  DFFQX1 \prev_key1_reg_reg[70]  ( .D(n3842), .CK(clk), .Q(prev_key1_reg[70])
         );
  DFFQX1 \prev_key1_reg_reg[69]  ( .D(n3843), .CK(clk), .Q(prev_key1_reg[69])
         );
  DFFQX1 \prev_key1_reg_reg[67]  ( .D(n3845), .CK(clk), .Q(prev_key1_reg[67])
         );
  DFFQX1 \prev_key1_reg_reg[66]  ( .D(n3846), .CK(clk), .Q(prev_key1_reg[66])
         );
  DFFRX1 ready_reg_reg ( .D(n1737), .CK(clk), .RN(n4407), .Q(ready) );
  DFFRX1 \key_mem_reg[3][107]  ( .D(n2142), .CK(clk), .RN(n4471), .Q(
        \key_mem[3][107] ) );
  DFFRX1 \key_mem_reg[7][107]  ( .D(n2654), .CK(clk), .RN(n4470), .Q(
        \key_mem[7][107] ) );
  DFFRX1 \key_mem_reg[11][107]  ( .D(n3166), .CK(clk), .RN(n4479), .Q(
        \key_mem[11][107] ) );
  DFFRX1 \key_mem_reg[3][19]  ( .D(n2230), .CK(clk), .RN(n4426), .Q(
        \key_mem[3][19] ) );
  DFFRX1 \key_mem_reg[7][19]  ( .D(n2742), .CK(clk), .RN(n4446), .Q(
        \key_mem[7][19] ) );
  DFFRX1 \key_mem_reg[11][19]  ( .D(n3254), .CK(clk), .RN(n4443), .Q(
        \key_mem[11][19] ) );
  DFFRX1 \key_mem_reg[2][107]  ( .D(n2014), .CK(clk), .RN(n4466), .Q(
        \key_mem[2][107] ) );
  DFFRX1 \key_mem_reg[6][107]  ( .D(n2526), .CK(clk), .RN(n4564), .Q(
        \key_mem[6][107] ) );
  DFFRX1 \key_mem_reg[10][107]  ( .D(n3038), .CK(clk), .RN(n4478), .Q(
        \key_mem[10][107] ) );
  DFFRX1 \key_mem_reg[2][19]  ( .D(n2102), .CK(clk), .RN(n4423), .Q(
        \key_mem[2][19] ) );
  DFFRX1 \key_mem_reg[6][19]  ( .D(n2614), .CK(clk), .RN(n4444), .Q(
        \key_mem[6][19] ) );
  DFFRX1 \key_mem_reg[10][19]  ( .D(n3126), .CK(clk), .RN(n4441), .Q(
        \key_mem[10][19] ) );
  DFFRX1 \key_mem_reg[13][107]  ( .D(n3422), .CK(clk), .RN(n4477), .Q(
        \key_mem[13][107] ) );
  DFFRX1 \key_mem_reg[13][19]  ( .D(n3510), .CK(clk), .RN(n4554), .Q(
        \key_mem[13][19] ) );
  DFFRX1 \key_mem_reg[12][107]  ( .D(n3294), .CK(clk), .RN(n4476), .Q(
        \key_mem[12][107] ) );
  DFFRX1 \key_mem_reg[12][19]  ( .D(n3382), .CK(clk), .RN(n4483), .Q(
        \key_mem[12][19] ) );
  DFFX1 \prev_key0_reg_reg[87]  ( .D(n3697), .CK(clk), .QN(n171) );
  DFFX1 \prev_key0_reg_reg[86]  ( .D(n3698), .CK(clk), .QN(n172) );
  DFFX1 \prev_key0_reg_reg[85]  ( .D(n3699), .CK(clk), .QN(n173) );
  DFFX1 \prev_key0_reg_reg[84]  ( .D(n3700), .CK(clk), .QN(n174) );
  DFFX1 \prev_key0_reg_reg[83]  ( .D(n3701), .CK(clk), .QN(n175) );
  DFFX1 \prev_key0_reg_reg[82]  ( .D(n3702), .CK(clk), .QN(n176) );
  DFFX1 \prev_key0_reg_reg[81]  ( .D(n3703), .CK(clk), .QN(n177) );
  DFFX1 \prev_key0_reg_reg[80]  ( .D(n3704), .CK(clk), .QN(n178) );
  DFFX1 \prev_key0_reg_reg[79]  ( .D(n3705), .CK(clk), .QN(n179) );
  DFFX1 \prev_key0_reg_reg[78]  ( .D(n3706), .CK(clk), .QN(n180) );
  DFFX1 \prev_key0_reg_reg[77]  ( .D(n3707), .CK(clk), .QN(n181) );
  DFFX1 \prev_key0_reg_reg[76]  ( .D(n3708), .CK(clk), .QN(n182) );
  DFFX1 \prev_key0_reg_reg[75]  ( .D(n3709), .CK(clk), .QN(n183) );
  DFFX1 \prev_key0_reg_reg[74]  ( .D(n3710), .CK(clk), .QN(n184) );
  DFFX1 \prev_key0_reg_reg[73]  ( .D(n3711), .CK(clk), .QN(n185) );
  DFFX1 \prev_key0_reg_reg[72]  ( .D(n3712), .CK(clk), .QN(n186) );
  DFFX1 \prev_key0_reg_reg[71]  ( .D(n3713), .CK(clk), .QN(n187) );
  DFFX1 \prev_key0_reg_reg[70]  ( .D(n3714), .CK(clk), .QN(n188) );
  DFFX1 \prev_key0_reg_reg[69]  ( .D(n3715), .CK(clk), .QN(n189) );
  DFFX1 \prev_key0_reg_reg[68]  ( .D(n3716), .CK(clk), .QN(n190) );
  DFFX1 \prev_key0_reg_reg[67]  ( .D(n3717), .CK(clk), .QN(n191) );
  DFFX1 \prev_key0_reg_reg[66]  ( .D(n3718), .CK(clk), .QN(n192) );
  DFFX1 \prev_key0_reg_reg[65]  ( .D(n3719), .CK(clk), .QN(n193) );
  DFFX1 \prev_key0_reg_reg[64]  ( .D(n3720), .CK(clk), .QN(n194) );
  DFFRX1 \rcon_reg_reg[1]  ( .D(n3919), .CK(clk), .RN(n4556), .QN(n293) );
  DFFRX1 \rcon_reg_reg[4]  ( .D(n3916), .CK(clk), .RN(n4471), .QN(n287) );
  DFFRX1 \rcon_reg_reg[5]  ( .D(n3915), .CK(clk), .RN(n4471), .QN(n285) );
  DFFRX1 \rcon_reg_reg[6]  ( .D(n3914), .CK(clk), .RN(n4471), .QN(n283) );
  DFFRX1 \rcon_reg_reg[7]  ( .D(n3921), .CK(clk), .RN(n4491), .Q(rcon_reg[7]), 
        .QN(n281) );
  DFFRX1 \rcon_reg_reg[2]  ( .D(n3918), .CK(clk), .RN(n4555), .Q(rcon_reg[2]), 
        .QN(n291) );
  DFFRX1 \rcon_reg_reg[3]  ( .D(n3917), .CK(clk), .RN(n4555), .Q(rcon_reg[3]), 
        .QN(n289) );
  DFFQX1 \prev_key0_reg_reg[23]  ( .D(n3761), .CK(clk), .Q(prev_key0_reg[23])
         );
  DFFQX1 \prev_key0_reg_reg[21]  ( .D(n3763), .CK(clk), .Q(prev_key0_reg[21])
         );
  DFFQX1 \prev_key0_reg_reg[19]  ( .D(n3765), .CK(clk), .Q(prev_key0_reg[19])
         );
  DFFQX1 \prev_key0_reg_reg[18]  ( .D(n3766), .CK(clk), .Q(prev_key0_reg[18])
         );
  DFFQX1 \prev_key0_reg_reg[15]  ( .D(n3769), .CK(clk), .Q(prev_key0_reg[15])
         );
  DFFQX1 \prev_key0_reg_reg[14]  ( .D(n3770), .CK(clk), .Q(prev_key0_reg[14])
         );
  DFFQX1 \prev_key0_reg_reg[13]  ( .D(n3771), .CK(clk), .Q(prev_key0_reg[13])
         );
  DFFQX1 \prev_key0_reg_reg[11]  ( .D(n3773), .CK(clk), .Q(prev_key0_reg[11])
         );
  DFFQX1 \prev_key0_reg_reg[10]  ( .D(n3774), .CK(clk), .Q(prev_key0_reg[10])
         );
  DFFQX1 \prev_key0_reg_reg[8]  ( .D(n3776), .CK(clk), .Q(prev_key0_reg[8]) );
  DFFQX1 \prev_key0_reg_reg[7]  ( .D(n3777), .CK(clk), .Q(prev_key0_reg[7]) );
  DFFQX1 \prev_key0_reg_reg[6]  ( .D(n3778), .CK(clk), .Q(prev_key0_reg[6]) );
  DFFQX1 \prev_key0_reg_reg[5]  ( .D(n3779), .CK(clk), .Q(prev_key0_reg[5]) );
  DFFQX1 \prev_key0_reg_reg[4]  ( .D(n3780), .CK(clk), .Q(prev_key0_reg[4]) );
  DFFQX1 \prev_key0_reg_reg[3]  ( .D(n3781), .CK(clk), .Q(prev_key0_reg[3]) );
  DFFQX1 \prev_key0_reg_reg[2]  ( .D(n3782), .CK(clk), .Q(prev_key0_reg[2]) );
  DFFQX1 \prev_key0_reg_reg[1]  ( .D(n3783), .CK(clk), .Q(prev_key0_reg[1]) );
  DFFQX1 \prev_key0_reg_reg[0]  ( .D(n3784), .CK(clk), .Q(prev_key0_reg[0]) );
  DFFQX1 \prev_key0_reg_reg[31]  ( .D(n3753), .CK(clk), .Q(prev_key0_reg[31])
         );
  DFFQX1 \prev_key0_reg_reg[24]  ( .D(n3760), .CK(clk), .Q(prev_key0_reg[24])
         );
  DFFQX1 \prev_key0_reg_reg[26]  ( .D(n3758), .CK(clk), .Q(prev_key0_reg[26])
         );
  DFFQX1 \prev_key0_reg_reg[27]  ( .D(n3757), .CK(clk), .Q(prev_key0_reg[27])
         );
  DFFQX1 \prev_key0_reg_reg[30]  ( .D(n3754), .CK(clk), .Q(prev_key0_reg[30])
         );
  DFFQX1 \prev_key0_reg_reg[29]  ( .D(n3755), .CK(clk), .Q(prev_key0_reg[29])
         );
  DFFQX1 \prev_key0_reg_reg[28]  ( .D(n3756), .CK(clk), .Q(prev_key0_reg[28])
         );
  DFFQX1 \prev_key0_reg_reg[25]  ( .D(n3759), .CK(clk), .Q(prev_key0_reg[25])
         );
  DFFQX1 \prev_key1_reg_reg[105]  ( .D(n3807), .CK(clk), .Q(prev_key1_reg[105]) );
  DFFQX1 \prev_key0_reg_reg[119]  ( .D(n3666), .CK(clk), .Q(prev_key0_reg[119]) );
  DFFQX1 \prev_key0_reg_reg[117]  ( .D(n3668), .CK(clk), .Q(prev_key0_reg[117]) );
  DFFQX1 \prev_key0_reg_reg[115]  ( .D(n3670), .CK(clk), .Q(prev_key0_reg[115]) );
  DFFQX1 \prev_key0_reg_reg[114]  ( .D(n3671), .CK(clk), .Q(prev_key0_reg[114]) );
  DFFQX1 \prev_key0_reg_reg[113]  ( .D(n3672), .CK(clk), .Q(prev_key0_reg[113]) );
  DFFQX1 \prev_key0_reg_reg[111]  ( .D(n3674), .CK(clk), .Q(prev_key0_reg[111]) );
  DFFQX1 \prev_key0_reg_reg[110]  ( .D(n3675), .CK(clk), .Q(prev_key0_reg[110]) );
  DFFQX1 \prev_key0_reg_reg[109]  ( .D(n3676), .CK(clk), .Q(prev_key0_reg[109]) );
  DFFQX1 \prev_key0_reg_reg[107]  ( .D(n3678), .CK(clk), .Q(prev_key0_reg[107]) );
  DFFQX1 \prev_key0_reg_reg[106]  ( .D(n3679), .CK(clk), .Q(prev_key0_reg[106]) );
  DFFQX1 \prev_key0_reg_reg[104]  ( .D(n3681), .CK(clk), .Q(prev_key0_reg[104]) );
  DFFQX1 \prev_key0_reg_reg[103]  ( .D(n3682), .CK(clk), .Q(prev_key0_reg[103]) );
  DFFQX1 \prev_key0_reg_reg[101]  ( .D(n3684), .CK(clk), .Q(prev_key0_reg[101]) );
  DFFQX1 \prev_key0_reg_reg[100]  ( .D(n3685), .CK(clk), .Q(prev_key0_reg[100]) );
  DFFQX1 \prev_key0_reg_reg[99]  ( .D(n3686), .CK(clk), .Q(prev_key0_reg[99])
         );
  DFFQX1 \prev_key0_reg_reg[98]  ( .D(n3913), .CK(clk), .Q(prev_key0_reg[98])
         );
  DFFQX1 \prev_key0_reg_reg[97]  ( .D(n3687), .CK(clk), .Q(prev_key0_reg[97])
         );
  DFFQX1 \prev_key0_reg_reg[96]  ( .D(n3688), .CK(clk), .Q(prev_key0_reg[96])
         );
  DFFQX1 \prev_key0_reg_reg[95]  ( .D(n3689), .CK(clk), .Q(prev_key0_reg[95])
         );
  DFFQX1 \prev_key0_reg_reg[88]  ( .D(n3696), .CK(clk), .Q(prev_key0_reg[88])
         );
  DFFQX1 \prev_key0_reg_reg[90]  ( .D(n3694), .CK(clk), .Q(prev_key0_reg[90])
         );
  DFFQX1 \prev_key0_reg_reg[91]  ( .D(n3693), .CK(clk), .Q(prev_key0_reg[91])
         );
  DFFQX1 \prev_key0_reg_reg[94]  ( .D(n3690), .CK(clk), .Q(prev_key0_reg[94])
         );
  DFFQX1 \prev_key0_reg_reg[93]  ( .D(n3691), .CK(clk), .Q(prev_key0_reg[93])
         );
  DFFQX1 \prev_key0_reg_reg[92]  ( .D(n3692), .CK(clk), .Q(prev_key0_reg[92])
         );
  DFFQX1 \prev_key0_reg_reg[89]  ( .D(n3695), .CK(clk), .Q(prev_key0_reg[89])
         );
  DFFQX1 \prev_key1_reg_reg[110]  ( .D(n3802), .CK(clk), .Q(prev_key1_reg[110]) );
  DFFQX1 \prev_key1_reg_reg[97]  ( .D(n3815), .CK(clk), .Q(prev_key1_reg[97])
         );
  DFFQX1 \prev_key1_reg_reg[119]  ( .D(n3793), .CK(clk), .Q(prev_key1_reg[119]) );
  DFFQX1 \prev_key1_reg_reg[117]  ( .D(n3795), .CK(clk), .Q(prev_key1_reg[117]) );
  DFFQX1 \prev_key1_reg_reg[116]  ( .D(n3796), .CK(clk), .Q(prev_key1_reg[116]) );
  DFFQX1 \prev_key1_reg_reg[115]  ( .D(n3797), .CK(clk), .Q(prev_key1_reg[115]) );
  DFFQX1 \prev_key1_reg_reg[114]  ( .D(n3798), .CK(clk), .Q(prev_key1_reg[114]) );
  DFFQX1 \prev_key1_reg_reg[113]  ( .D(n3799), .CK(clk), .Q(prev_key1_reg[113]) );
  DFFQX1 \prev_key1_reg_reg[112]  ( .D(n3800), .CK(clk), .Q(prev_key1_reg[112]) );
  DFFQX1 \prev_key1_reg_reg[111]  ( .D(n3801), .CK(clk), .Q(prev_key1_reg[111]) );
  DFFQX1 \prev_key1_reg_reg[109]  ( .D(n3803), .CK(clk), .Q(prev_key1_reg[109]) );
  DFFQX1 \prev_key1_reg_reg[107]  ( .D(n3805), .CK(clk), .Q(prev_key1_reg[107]) );
  DFFQX1 \prev_key1_reg_reg[106]  ( .D(n3806), .CK(clk), .Q(prev_key1_reg[106]) );
  DFFQX1 \prev_key1_reg_reg[104]  ( .D(n3808), .CK(clk), .Q(prev_key1_reg[104]) );
  DFFQX1 \prev_key1_reg_reg[103]  ( .D(n3809), .CK(clk), .Q(prev_key1_reg[103]) );
  DFFQX1 \prev_key1_reg_reg[102]  ( .D(n3810), .CK(clk), .Q(prev_key1_reg[102]) );
  DFFQX1 \prev_key1_reg_reg[101]  ( .D(n3811), .CK(clk), .Q(prev_key1_reg[101]) );
  DFFQX1 \prev_key1_reg_reg[100]  ( .D(n3812), .CK(clk), .Q(prev_key1_reg[100]) );
  DFFQX1 \prev_key1_reg_reg[99]  ( .D(n3813), .CK(clk), .Q(prev_key1_reg[99])
         );
  DFFQX1 \prev_key1_reg_reg[98]  ( .D(n3814), .CK(clk), .Q(prev_key1_reg[98])
         );
  DFFQX1 \prev_key1_reg_reg[96]  ( .D(n3816), .CK(clk), .Q(prev_key1_reg[96])
         );
  DFFQX1 \prev_key1_reg_reg[120]  ( .D(n3792), .CK(clk), .Q(prev_key1_reg[120]) );
  DFFQX1 \prev_key1_reg_reg[88]  ( .D(n3824), .CK(clk), .Q(prev_key1_reg[88])
         );
  DFFQX1 \prev_key1_reg_reg[122]  ( .D(n3790), .CK(clk), .Q(prev_key1_reg[122]) );
  DFFQX1 \prev_key1_reg_reg[90]  ( .D(n3822), .CK(clk), .Q(prev_key1_reg[90])
         );
  DFFQX1 \prev_key1_reg_reg[123]  ( .D(n3789), .CK(clk), .Q(prev_key1_reg[123]) );
  DFFQX1 \prev_key1_reg_reg[91]  ( .D(n3821), .CK(clk), .Q(prev_key1_reg[91])
         );
  DFFQX1 \prev_key1_reg_reg[126]  ( .D(n3786), .CK(clk), .Q(prev_key1_reg[126]) );
  DFFQX1 \prev_key1_reg_reg[94]  ( .D(n3818), .CK(clk), .Q(prev_key1_reg[94])
         );
  DFFQX1 \prev_key1_reg_reg[125]  ( .D(n3787), .CK(clk), .Q(prev_key1_reg[125]) );
  DFFQX1 \prev_key1_reg_reg[93]  ( .D(n3819), .CK(clk), .Q(prev_key1_reg[93])
         );
  DFFQX1 \prev_key1_reg_reg[124]  ( .D(n3788), .CK(clk), .Q(prev_key1_reg[124]) );
  DFFQX1 \prev_key1_reg_reg[92]  ( .D(n3820), .CK(clk), .Q(prev_key1_reg[92])
         );
  DFFQX1 \prev_key1_reg_reg[121]  ( .D(n3791), .CK(clk), .Q(prev_key1_reg[121]) );
  DFFQX1 \prev_key1_reg_reg[89]  ( .D(n3823), .CK(clk), .Q(prev_key1_reg[89])
         );
  DFFQX1 \prev_key0_reg_reg[127]  ( .D(n3658), .CK(clk), .Q(prev_key0_reg[127]) );
  DFFQX1 \prev_key0_reg_reg[120]  ( .D(n3665), .CK(clk), .Q(prev_key0_reg[120]) );
  DFFQX1 \prev_key0_reg_reg[122]  ( .D(n3663), .CK(clk), .Q(prev_key0_reg[122]) );
  DFFQX1 \prev_key0_reg_reg[123]  ( .D(n3662), .CK(clk), .Q(prev_key0_reg[123]) );
  DFFQX1 \prev_key0_reg_reg[126]  ( .D(n3659), .CK(clk), .Q(prev_key0_reg[126]) );
  DFFQX1 \prev_key0_reg_reg[125]  ( .D(n3660), .CK(clk), .Q(prev_key0_reg[125]) );
  DFFQX1 \prev_key0_reg_reg[124]  ( .D(n3661), .CK(clk), .Q(prev_key0_reg[124]) );
  DFFQX1 \prev_key0_reg_reg[121]  ( .D(n3664), .CK(clk), .Q(prev_key0_reg[121]) );
  DFFQX1 \prev_key0_reg_reg[55]  ( .D(n3729), .CK(clk), .Q(prev_key0_reg[55])
         );
  DFFQX1 \prev_key0_reg_reg[53]  ( .D(n3731), .CK(clk), .Q(prev_key0_reg[53])
         );
  DFFQX1 \prev_key0_reg_reg[51]  ( .D(n3733), .CK(clk), .Q(prev_key0_reg[51])
         );
  DFFQX1 \prev_key0_reg_reg[50]  ( .D(n3734), .CK(clk), .Q(prev_key0_reg[50])
         );
  DFFQX1 \prev_key0_reg_reg[47]  ( .D(n3737), .CK(clk), .Q(prev_key0_reg[47])
         );
  DFFQX1 \prev_key0_reg_reg[46]  ( .D(n3738), .CK(clk), .Q(prev_key0_reg[46])
         );
  DFFQX1 \prev_key0_reg_reg[45]  ( .D(n3739), .CK(clk), .Q(prev_key0_reg[45])
         );
  DFFQX1 \prev_key0_reg_reg[43]  ( .D(n3741), .CK(clk), .Q(prev_key0_reg[43])
         );
  DFFQX1 \prev_key0_reg_reg[42]  ( .D(n3742), .CK(clk), .Q(prev_key0_reg[42])
         );
  DFFQX1 \prev_key0_reg_reg[56]  ( .D(n3728), .CK(clk), .Q(prev_key0_reg[56])
         );
  DFFQX1 \prev_key0_reg_reg[58]  ( .D(n3726), .CK(clk), .Q(prev_key0_reg[58])
         );
  DFFQX1 \prev_key0_reg_reg[59]  ( .D(n3725), .CK(clk), .Q(prev_key0_reg[59])
         );
  DFFQX1 \prev_key0_reg_reg[62]  ( .D(n3722), .CK(clk), .Q(prev_key0_reg[62])
         );
  DFFQX1 \prev_key0_reg_reg[61]  ( .D(n3723), .CK(clk), .Q(prev_key0_reg[61])
         );
  DFFQX1 \prev_key0_reg_reg[60]  ( .D(n3724), .CK(clk), .Q(prev_key0_reg[60])
         );
  DFFQX1 \prev_key0_reg_reg[57]  ( .D(n3727), .CK(clk), .Q(prev_key0_reg[57])
         );
  DFFQX1 \prev_key0_reg_reg[102]  ( .D(n3683), .CK(clk), .Q(prev_key0_reg[102]) );
  DFFRX1 \rcon_reg_reg[0]  ( .D(n3920), .CK(clk), .RN(n4461), .QN(n295) );
  DFFRX1 \key_mem_reg[5][119]  ( .D(n2386), .CK(clk), .RN(n4430), .Q(
        \key_mem[5][119] ) );
  DFFRX1 \key_mem_reg[9][119]  ( .D(n2898), .CK(clk), .RN(n4431), .Q(
        \key_mem[9][119] ) );
  DFFRX1 \key_mem_reg[5][118]  ( .D(n2387), .CK(clk), .RN(n4432), .Q(
        \key_mem[5][118] ) );
  DFFRX1 \key_mem_reg[9][118]  ( .D(n2899), .CK(clk), .RN(n4432), .Q(
        \key_mem[9][118] ) );
  DFFRX1 \key_mem_reg[5][117]  ( .D(n2388), .CK(clk), .RN(n4433), .Q(
        \key_mem[5][117] ) );
  DFFRX1 \key_mem_reg[9][117]  ( .D(n2900), .CK(clk), .RN(n4433), .Q(
        \key_mem[9][117] ) );
  DFFRX1 \key_mem_reg[5][116]  ( .D(n2389), .CK(clk), .RN(n4499), .Q(
        \key_mem[5][116] ) );
  DFFRX1 \key_mem_reg[9][116]  ( .D(n2901), .CK(clk), .RN(n4405), .Q(
        \key_mem[9][116] ) );
  DFFRX1 \key_mem_reg[5][115]  ( .D(n2390), .CK(clk), .RN(n4397), .Q(
        \key_mem[5][115] ) );
  DFFRX1 \key_mem_reg[9][115]  ( .D(n2902), .CK(clk), .RN(n4434), .Q(
        \key_mem[9][115] ) );
  DFFRX1 \key_mem_reg[5][114]  ( .D(n2391), .CK(clk), .RN(n4435), .Q(
        \key_mem[5][114] ) );
  DFFRX1 \key_mem_reg[9][114]  ( .D(n2903), .CK(clk), .RN(n4436), .Q(
        \key_mem[9][114] ) );
  DFFRX1 \key_mem_reg[5][113]  ( .D(n2392), .CK(clk), .RN(n4437), .Q(
        \key_mem[5][113] ) );
  DFFRX1 \key_mem_reg[9][113]  ( .D(n2904), .CK(clk), .RN(n4437), .Q(
        \key_mem[9][113] ) );
  DFFRX1 \key_mem_reg[5][112]  ( .D(n2393), .CK(clk), .RN(n4439), .Q(
        \key_mem[5][112] ) );
  DFFRX1 \key_mem_reg[9][112]  ( .D(n2905), .CK(clk), .RN(n4439), .Q(
        \key_mem[9][112] ) );
  DFFRX1 \key_mem_reg[5][111]  ( .D(n2394), .CK(clk), .RN(n4475), .Q(
        \key_mem[5][111] ) );
  DFFRX1 \key_mem_reg[9][111]  ( .D(n2906), .CK(clk), .RN(n4418), .Q(
        \key_mem[9][111] ) );
  DFFRX1 \key_mem_reg[5][110]  ( .D(n2395), .CK(clk), .RN(n4442), .Q(
        \key_mem[5][110] ) );
  DFFRX1 \key_mem_reg[9][110]  ( .D(n2907), .CK(clk), .RN(n4439), .Q(
        \key_mem[9][110] ) );
  DFFRX1 \key_mem_reg[5][109]  ( .D(n2396), .CK(clk), .RN(n4420), .Q(
        \key_mem[5][109] ) );
  DFFRX1 \key_mem_reg[9][109]  ( .D(n2908), .CK(clk), .RN(n4420), .Q(
        \key_mem[9][109] ) );
  DFFRX1 \key_mem_reg[5][108]  ( .D(n2397), .CK(clk), .RN(n4421), .Q(
        \key_mem[5][108] ) );
  DFFRX1 \key_mem_reg[9][108]  ( .D(n2909), .CK(clk), .RN(n4422), .Q(
        \key_mem[9][108] ) );
  DFFRX1 \key_mem_reg[5][107]  ( .D(n2398), .CK(clk), .RN(n4464), .Q(
        \key_mem[5][107] ) );
  DFFRX1 \key_mem_reg[9][107]  ( .D(n2910), .CK(clk), .RN(n4474), .Q(
        \key_mem[9][107] ) );
  DFFRX1 \key_mem_reg[5][106]  ( .D(n2399), .CK(clk), .RN(n4423), .Q(
        \key_mem[5][106] ) );
  DFFRX1 \key_mem_reg[9][106]  ( .D(n2911), .CK(clk), .RN(n4423), .Q(
        \key_mem[9][106] ) );
  DFFRX1 \key_mem_reg[5][105]  ( .D(n2400), .CK(clk), .RN(n4425), .Q(
        \key_mem[5][105] ) );
  DFFRX1 \key_mem_reg[9][105]  ( .D(n2912), .CK(clk), .RN(n4425), .Q(
        \key_mem[9][105] ) );
  DFFRX1 \key_mem_reg[5][104]  ( .D(n2401), .CK(clk), .RN(n4426), .Q(
        \key_mem[5][104] ) );
  DFFRX1 \key_mem_reg[9][104]  ( .D(n2913), .CK(clk), .RN(n4427), .Q(
        \key_mem[9][104] ) );
  DFFRX1 \key_mem_reg[5][103]  ( .D(n2402), .CK(clk), .RN(n4428), .Q(
        \key_mem[5][103] ) );
  DFFRX1 \key_mem_reg[9][103]  ( .D(n2914), .CK(clk), .RN(n4429), .Q(
        \key_mem[9][103] ) );
  DFFRX1 \key_mem_reg[5][102]  ( .D(n2403), .CK(clk), .RN(n4456), .Q(
        \key_mem[5][102] ) );
  DFFRX1 \key_mem_reg[9][102]  ( .D(n2915), .CK(clk), .RN(n4457), .Q(
        \key_mem[9][102] ) );
  DFFRX1 \key_mem_reg[5][101]  ( .D(n2404), .CK(clk), .RN(n4458), .Q(
        \key_mem[5][101] ) );
  DFFRX1 \key_mem_reg[9][101]  ( .D(n2916), .CK(clk), .RN(n4458), .Q(
        \key_mem[9][101] ) );
  DFFRX1 \key_mem_reg[5][100]  ( .D(n2405), .CK(clk), .RN(n4460), .Q(
        \key_mem[5][100] ) );
  DFFRX1 \key_mem_reg[9][100]  ( .D(n2917), .CK(clk), .RN(n4460), .Q(
        \key_mem[9][100] ) );
  DFFRX1 \key_mem_reg[5][99]  ( .D(n2406), .CK(clk), .RN(n4469), .Q(
        \key_mem[5][99] ) );
  DFFRX1 \key_mem_reg[9][99]  ( .D(n2918), .CK(clk), .RN(n4461), .Q(
        \key_mem[9][99] ) );
  DFFRX1 \key_mem_reg[5][98]  ( .D(n2407), .CK(clk), .RN(n4462), .Q(
        \key_mem[5][98] ) );
  DFFRX1 \key_mem_reg[9][98]  ( .D(n2919), .CK(clk), .RN(n4463), .Q(
        \key_mem[9][98] ) );
  DFFRX1 \key_mem_reg[5][97]  ( .D(n2408), .CK(clk), .RN(n4464), .Q(
        \key_mem[5][97] ) );
  DFFRX1 \key_mem_reg[9][97]  ( .D(n2920), .CK(clk), .RN(n4464), .Q(
        \key_mem[9][97] ) );
  DFFRX1 \key_mem_reg[5][96]  ( .D(n2409), .CK(clk), .RN(n4466), .Q(
        \key_mem[5][96] ) );
  DFFRX1 \key_mem_reg[9][96]  ( .D(n2921), .CK(clk), .RN(n4466), .Q(
        \key_mem[9][96] ) );
  DFFRX1 \key_mem_reg[5][87]  ( .D(n2418), .CK(clk), .RN(n4467), .Q(
        \key_mem[5][87] ) );
  DFFRX1 \key_mem_reg[9][87]  ( .D(n2930), .CK(clk), .RN(n4468), .Q(
        \key_mem[9][87] ) );
  DFFRX1 \key_mem_reg[5][86]  ( .D(n2419), .CK(clk), .RN(n4469), .Q(
        \key_mem[5][86] ) );
  DFFRX1 \key_mem_reg[9][86]  ( .D(n2931), .CK(clk), .RN(n4440), .Q(
        \key_mem[9][86] ) );
  DFFRX1 \key_mem_reg[5][85]  ( .D(n2420), .CK(clk), .RN(n4442), .Q(
        \key_mem[5][85] ) );
  DFFRX1 \key_mem_reg[9][85]  ( .D(n2932), .CK(clk), .RN(n4442), .Q(
        \key_mem[9][85] ) );
  DFFRX1 \key_mem_reg[5][84]  ( .D(n2421), .CK(clk), .RN(n4443), .Q(
        \key_mem[5][84] ) );
  DFFRX1 \key_mem_reg[9][84]  ( .D(n2933), .CK(clk), .RN(n4444), .Q(
        \key_mem[9][84] ) );
  DFFRX1 \key_mem_reg[5][83]  ( .D(n2422), .CK(clk), .RN(n4445), .Q(
        \key_mem[5][83] ) );
  DFFRX1 \key_mem_reg[9][83]  ( .D(n2934), .CK(clk), .RN(n4446), .Q(
        \key_mem[9][83] ) );
  DFFRX1 \key_mem_reg[5][82]  ( .D(n2423), .CK(clk), .RN(n4447), .Q(
        \key_mem[5][82] ) );
  DFFRX1 \key_mem_reg[9][82]  ( .D(n2935), .CK(clk), .RN(n4447), .Q(
        \key_mem[9][82] ) );
  DFFRX1 \key_mem_reg[5][81]  ( .D(n2424), .CK(clk), .RN(n4449), .Q(
        \key_mem[5][81] ) );
  DFFRX1 \key_mem_reg[9][81]  ( .D(n2936), .CK(clk), .RN(n4449), .Q(
        \key_mem[9][81] ) );
  DFFRX1 \key_mem_reg[5][80]  ( .D(n2425), .CK(clk), .RN(n4451), .Q(
        \key_mem[5][80] ) );
  DFFRX1 \key_mem_reg[9][80]  ( .D(n2937), .CK(clk), .RN(n4451), .Q(
        \key_mem[9][80] ) );
  DFFRX1 \key_mem_reg[5][79]  ( .D(n2426), .CK(clk), .RN(n4452), .Q(
        \key_mem[5][79] ) );
  DFFRX1 \key_mem_reg[9][79]  ( .D(n2938), .CK(clk), .RN(n4453), .Q(
        \key_mem[9][79] ) );
  DFFRX1 \key_mem_reg[5][78]  ( .D(n2427), .CK(clk), .RN(n4454), .Q(
        \key_mem[5][78] ) );
  DFFRX1 \key_mem_reg[9][78]  ( .D(n2939), .CK(clk), .RN(n4455), .Q(
        \key_mem[9][78] ) );
  DFFRX1 \key_mem_reg[5][77]  ( .D(n2428), .CK(clk), .RN(n4373), .Q(
        \key_mem[5][77] ) );
  DFFRX1 \key_mem_reg[9][77]  ( .D(n2940), .CK(clk), .RN(n4373), .Q(
        \key_mem[9][77] ) );
  DFFRX1 \key_mem_reg[5][76]  ( .D(n2429), .CK(clk), .RN(n4375), .Q(
        \key_mem[5][76] ) );
  DFFRX1 \key_mem_reg[9][76]  ( .D(n2941), .CK(clk), .RN(n4375), .Q(
        \key_mem[9][76] ) );
  DFFRX1 \key_mem_reg[5][75]  ( .D(n2430), .CK(clk), .RN(n4376), .Q(
        \key_mem[5][75] ) );
  DFFRX1 \key_mem_reg[9][75]  ( .D(n2942), .CK(clk), .RN(n4377), .Q(
        \key_mem[9][75] ) );
  DFFRX1 \key_mem_reg[5][74]  ( .D(n2431), .CK(clk), .RN(n4378), .Q(
        \key_mem[5][74] ) );
  DFFRX1 \key_mem_reg[9][74]  ( .D(n2943), .CK(clk), .RN(n4379), .Q(
        \key_mem[9][74] ) );
  DFFRX1 \key_mem_reg[5][73]  ( .D(n2432), .CK(clk), .RN(n4380), .Q(
        \key_mem[5][73] ) );
  DFFRX1 \key_mem_reg[9][73]  ( .D(n2944), .CK(clk), .RN(n4380), .Q(
        \key_mem[9][73] ) );
  DFFRX1 \key_mem_reg[5][72]  ( .D(n2433), .CK(clk), .RN(n4382), .Q(
        \key_mem[5][72] ) );
  DFFRX1 \key_mem_reg[9][72]  ( .D(n2945), .CK(clk), .RN(n4382), .Q(
        \key_mem[9][72] ) );
  DFFRX1 \key_mem_reg[5][71]  ( .D(n2434), .CK(clk), .RN(n4383), .Q(
        \key_mem[5][71] ) );
  DFFRX1 \key_mem_reg[9][71]  ( .D(n2946), .CK(clk), .RN(n4384), .Q(
        \key_mem[9][71] ) );
  DFFRX1 \key_mem_reg[5][70]  ( .D(n2435), .CK(clk), .RN(n4385), .Q(
        \key_mem[5][70] ) );
  DFFRX1 \key_mem_reg[9][70]  ( .D(n2947), .CK(clk), .RN(n4386), .Q(
        \key_mem[9][70] ) );
  DFFRX1 \key_mem_reg[5][69]  ( .D(n2436), .CK(clk), .RN(n4387), .Q(
        \key_mem[5][69] ) );
  DFFRX1 \key_mem_reg[9][69]  ( .D(n2948), .CK(clk), .RN(n4387), .Q(
        \key_mem[9][69] ) );
  DFFRX1 \key_mem_reg[5][68]  ( .D(n2437), .CK(clk), .RN(n4408), .Q(
        \key_mem[5][68] ) );
  DFFRX1 \key_mem_reg[9][68]  ( .D(n2949), .CK(clk), .RN(n4459), .Q(
        \key_mem[9][68] ) );
  DFFRX1 \key_mem_reg[5][67]  ( .D(n2438), .CK(clk), .RN(n4559), .Q(
        \key_mem[5][67] ) );
  DFFRX1 \key_mem_reg[9][67]  ( .D(n2950), .CK(clk), .RN(n4380), .Q(
        \key_mem[9][67] ) );
  DFFRX1 \key_mem_reg[5][66]  ( .D(n2439), .CK(clk), .RN(n4400), .Q(
        \key_mem[5][66] ) );
  DFFRX1 \key_mem_reg[9][66]  ( .D(n2951), .CK(clk), .RN(n4390), .Q(
        \key_mem[9][66] ) );
  DFFRX1 \key_mem_reg[5][65]  ( .D(n2440), .CK(clk), .RN(n4457), .Q(
        \key_mem[5][65] ) );
  DFFRX1 \key_mem_reg[9][65]  ( .D(n2952), .CK(clk), .RN(n4458), .Q(
        \key_mem[9][65] ) );
  DFFRX1 \key_mem_reg[5][64]  ( .D(n2441), .CK(clk), .RN(n4424), .Q(
        \key_mem[5][64] ) );
  DFFRX1 \key_mem_reg[9][64]  ( .D(n2953), .CK(clk), .RN(n4421), .Q(
        \key_mem[9][64] ) );
  DFFRX1 \key_mem_reg[5][55]  ( .D(n2450), .CK(clk), .RN(n4504), .Q(
        \key_mem[5][55] ) );
  DFFRX1 \key_mem_reg[9][55]  ( .D(n2962), .CK(clk), .RN(n4548), .Q(
        \key_mem[9][55] ) );
  DFFRX1 \key_mem_reg[5][54]  ( .D(n2451), .CK(clk), .RN(n4543), .Q(
        \key_mem[5][54] ) );
  DFFRX1 \key_mem_reg[9][54]  ( .D(n2963), .CK(clk), .RN(n4370), .Q(
        \key_mem[9][54] ) );
  DFFRX1 \key_mem_reg[5][53]  ( .D(n2452), .CK(clk), .RN(n4371), .Q(
        \key_mem[5][53] ) );
  DFFRX1 \key_mem_reg[9][53]  ( .D(n2964), .CK(clk), .RN(n4371), .Q(
        \key_mem[9][53] ) );
  DFFRX1 \key_mem_reg[5][52]  ( .D(n2453), .CK(clk), .RN(n4373), .Q(
        \key_mem[5][52] ) );
  DFFRX1 \key_mem_reg[9][52]  ( .D(n2965), .CK(clk), .RN(n4403), .Q(
        \key_mem[9][52] ) );
  DFFRX1 \key_mem_reg[5][51]  ( .D(n2454), .CK(clk), .RN(n4405), .Q(
        \key_mem[5][51] ) );
  DFFRX1 \key_mem_reg[9][51]  ( .D(n2966), .CK(clk), .RN(n4405), .Q(
        \key_mem[9][51] ) );
  DFFRX1 \key_mem_reg[5][50]  ( .D(n2455), .CK(clk), .RN(n4406), .Q(
        \key_mem[5][50] ) );
  DFFRX1 \key_mem_reg[9][50]  ( .D(n2967), .CK(clk), .RN(n4407), .Q(
        \key_mem[9][50] ) );
  DFFRX1 \key_mem_reg[5][49]  ( .D(n2456), .CK(clk), .RN(n4408), .Q(
        \key_mem[5][49] ) );
  DFFRX1 \key_mem_reg[9][49]  ( .D(n2968), .CK(clk), .RN(n4409), .Q(
        \key_mem[9][49] ) );
  DFFRX1 \key_mem_reg[5][47]  ( .D(n2458), .CK(clk), .RN(n4412), .Q(
        \key_mem[5][47] ) );
  DFFRX1 \key_mem_reg[9][47]  ( .D(n2970), .CK(clk), .RN(n4412), .Q(
        \key_mem[9][47] ) );
  DFFRX1 \key_mem_reg[5][46]  ( .D(n2459), .CK(clk), .RN(n4413), .Q(
        \key_mem[5][46] ) );
  DFFRX1 \key_mem_reg[9][46]  ( .D(n2971), .CK(clk), .RN(n4412), .Q(
        \key_mem[9][46] ) );
  DFFRX1 \key_mem_reg[5][45]  ( .D(n2460), .CK(clk), .RN(n4414), .Q(
        \key_mem[5][45] ) );
  DFFRX1 \key_mem_reg[9][45]  ( .D(n2972), .CK(clk), .RN(n4415), .Q(
        \key_mem[9][45] ) );
  DFFRX1 \key_mem_reg[5][44]  ( .D(n2461), .CK(clk), .RN(n4416), .Q(
        \key_mem[5][44] ) );
  DFFRX1 \key_mem_reg[9][44]  ( .D(n2973), .CK(clk), .RN(n4416), .Q(
        \key_mem[9][44] ) );
  DFFRX1 \key_mem_reg[5][43]  ( .D(n2462), .CK(clk), .RN(n4388), .Q(
        \key_mem[5][43] ) );
  DFFRX1 \key_mem_reg[9][43]  ( .D(n2974), .CK(clk), .RN(n4389), .Q(
        \key_mem[9][43] ) );
  DFFRX1 \key_mem_reg[5][42]  ( .D(n2463), .CK(clk), .RN(n4390), .Q(
        \key_mem[5][42] ) );
  DFFRX1 \key_mem_reg[9][42]  ( .D(n2975), .CK(clk), .RN(n4391), .Q(
        \key_mem[9][42] ) );
  DFFRX1 \key_mem_reg[5][41]  ( .D(n2464), .CK(clk), .RN(n4392), .Q(
        \key_mem[5][41] ) );
  DFFRX1 \key_mem_reg[9][41]  ( .D(n2976), .CK(clk), .RN(n4392), .Q(
        \key_mem[9][41] ) );
  DFFRX1 \key_mem_reg[5][40]  ( .D(n2465), .CK(clk), .RN(n4394), .Q(
        \key_mem[5][40] ) );
  DFFRX1 \key_mem_reg[9][40]  ( .D(n2977), .CK(clk), .RN(n4394), .Q(
        \key_mem[9][40] ) );
  DFFRX1 \key_mem_reg[5][39]  ( .D(n2466), .CK(clk), .RN(n4396), .Q(
        \key_mem[5][39] ) );
  DFFRX1 \key_mem_reg[9][39]  ( .D(n2978), .CK(clk), .RN(n4396), .Q(
        \key_mem[9][39] ) );
  DFFRX1 \key_mem_reg[5][38]  ( .D(n2467), .CK(clk), .RN(n4397), .Q(
        \key_mem[5][38] ) );
  DFFRX1 \key_mem_reg[9][38]  ( .D(n2979), .CK(clk), .RN(n4398), .Q(
        \key_mem[9][38] ) );
  DFFRX1 \key_mem_reg[5][37]  ( .D(n2468), .CK(clk), .RN(n4399), .Q(
        \key_mem[5][37] ) );
  DFFRX1 \key_mem_reg[9][37]  ( .D(n2980), .CK(clk), .RN(n4400), .Q(
        \key_mem[9][37] ) );
  DFFRX1 \key_mem_reg[5][36]  ( .D(n2469), .CK(clk), .RN(n4401), .Q(
        \key_mem[5][36] ) );
  DFFRX1 \key_mem_reg[9][36]  ( .D(n2981), .CK(clk), .RN(n4401), .Q(
        \key_mem[9][36] ) );
  DFFRX1 \key_mem_reg[5][35]  ( .D(n2470), .CK(clk), .RN(n4403), .Q(
        \key_mem[5][35] ) );
  DFFRX1 \key_mem_reg[9][35]  ( .D(n2982), .CK(clk), .RN(n4417), .Q(
        \key_mem[9][35] ) );
  DFFRX1 \key_mem_reg[5][34]  ( .D(n2471), .CK(clk), .RN(n4542), .Q(
        \key_mem[5][34] ) );
  DFFRX1 \key_mem_reg[9][34]  ( .D(n2983), .CK(clk), .RN(n4543), .Q(
        \key_mem[9][34] ) );
  DFFRX1 \key_mem_reg[5][33]  ( .D(n2472), .CK(clk), .RN(n4544), .Q(
        \key_mem[5][33] ) );
  DFFRX1 \key_mem_reg[9][33]  ( .D(n2984), .CK(clk), .RN(n4544), .Q(
        \key_mem[9][33] ) );
  DFFRX1 \key_mem_reg[5][32]  ( .D(n2473), .CK(clk), .RN(n4546), .Q(
        \key_mem[5][32] ) );
  DFFRX1 \key_mem_reg[9][32]  ( .D(n2985), .CK(clk), .RN(n4546), .Q(
        \key_mem[9][32] ) );
  DFFRX1 \key_mem_reg[5][23]  ( .D(n2482), .CK(clk), .RN(n4547), .Q(
        \key_mem[5][23] ) );
  DFFRX1 \key_mem_reg[9][23]  ( .D(n2994), .CK(clk), .RN(n4548), .Q(
        \key_mem[9][23] ) );
  DFFRX1 \key_mem_reg[5][22]  ( .D(n2483), .CK(clk), .RN(n4549), .Q(
        \key_mem[5][22] ) );
  DFFRX1 \key_mem_reg[9][22]  ( .D(n2995), .CK(clk), .RN(n4550), .Q(
        \key_mem[9][22] ) );
  DFFRX1 \key_mem_reg[5][21]  ( .D(n2484), .CK(clk), .RN(n4551), .Q(
        \key_mem[5][21] ) );
  DFFRX1 \key_mem_reg[9][21]  ( .D(n2996), .CK(clk), .RN(n4552), .Q(
        \key_mem[9][21] ) );
  DFFRX1 \key_mem_reg[5][20]  ( .D(n2485), .CK(clk), .RN(n4553), .Q(
        \key_mem[5][20] ) );
  DFFRX1 \key_mem_reg[9][20]  ( .D(n2997), .CK(clk), .RN(n4553), .Q(
        \key_mem[9][20] ) );
  DFFRX1 \key_mem_reg[5][19]  ( .D(n2486), .CK(clk), .RN(n4482), .Q(
        \key_mem[5][19] ) );
  DFFRX1 \key_mem_reg[9][19]  ( .D(n2998), .CK(clk), .RN(n4481), .Q(
        \key_mem[9][19] ) );
  DFFRX1 \key_mem_reg[5][18]  ( .D(n2487), .CK(clk), .RN(n4534), .Q(
        \key_mem[5][18] ) );
  DFFRX1 \key_mem_reg[9][18]  ( .D(n2999), .CK(clk), .RN(n4527), .Q(
        \key_mem[9][18] ) );
  DFFRX1 \key_mem_reg[5][16]  ( .D(n2489), .CK(clk), .RN(n4530), .Q(
        \key_mem[5][16] ) );
  DFFRX1 \key_mem_reg[9][16]  ( .D(n3001), .CK(clk), .RN(n4530), .Q(
        \key_mem[9][16] ) );
  DFFRX1 \key_mem_reg[5][15]  ( .D(n2490), .CK(clk), .RN(n4531), .Q(
        \key_mem[5][15] ) );
  DFFRX1 \key_mem_reg[9][15]  ( .D(n3002), .CK(clk), .RN(n4532), .Q(
        \key_mem[9][15] ) );
  DFFRX1 \key_mem_reg[5][14]  ( .D(n2491), .CK(clk), .RN(n4533), .Q(
        \key_mem[5][14] ) );
  DFFRX1 \key_mem_reg[9][14]  ( .D(n3003), .CK(clk), .RN(n4534), .Q(
        \key_mem[9][14] ) );
  DFFRX1 \key_mem_reg[5][13]  ( .D(n2492), .CK(clk), .RN(n4535), .Q(
        \key_mem[5][13] ) );
  DFFRX1 \key_mem_reg[9][13]  ( .D(n3004), .CK(clk), .RN(n4535), .Q(
        \key_mem[9][13] ) );
  DFFRX1 \key_mem_reg[5][12]  ( .D(n2493), .CK(clk), .RN(n4537), .Q(
        \key_mem[5][12] ) );
  DFFRX1 \key_mem_reg[9][12]  ( .D(n3005), .CK(clk), .RN(n4537), .Q(
        \key_mem[9][12] ) );
  DFFRX1 \key_mem_reg[5][11]  ( .D(n2494), .CK(clk), .RN(n4538), .Q(
        \key_mem[5][11] ) );
  DFFRX1 \key_mem_reg[9][11]  ( .D(n3006), .CK(clk), .RN(n4539), .Q(
        \key_mem[9][11] ) );
  DFFRX1 \key_mem_reg[5][10]  ( .D(n2495), .CK(clk), .RN(n4540), .Q(
        \key_mem[5][10] ) );
  DFFRX1 \key_mem_reg[9][10]  ( .D(n3007), .CK(clk), .RN(n4541), .Q(
        \key_mem[9][10] ) );
  DFFRX1 \key_mem_reg[5][9]  ( .D(n2496), .CK(clk), .RN(n4537), .Q(
        \key_mem[5][9] ) );
  DFFRX1 \key_mem_reg[9][9]  ( .D(n3008), .CK(clk), .RN(n4531), .Q(
        \key_mem[9][9] ) );
  DFFRX1 \key_mem_reg[5][8]  ( .D(n2497), .CK(clk), .RN(n4498), .Q(
        \key_mem[5][8] ) );
  DFFRX1 \key_mem_reg[9][8]  ( .D(n3009), .CK(clk), .RN(n4522), .Q(
        \key_mem[9][8] ) );
  DFFRX1 \key_mem_reg[5][7]  ( .D(n2498), .CK(clk), .RN(n4560), .Q(
        \key_mem[5][7] ) );
  DFFRX1 \key_mem_reg[9][7]  ( .D(n3010), .CK(clk), .RN(n4560), .Q(
        \key_mem[9][7] ) );
  DFFRX1 \key_mem_reg[5][6]  ( .D(n2499), .CK(clk), .RN(n4561), .Q(
        \key_mem[5][6] ) );
  DFFRX1 \key_mem_reg[9][6]  ( .D(n3011), .CK(clk), .RN(n4562), .Q(
        \key_mem[9][6] ) );
  DFFRX1 \key_mem_reg[5][5]  ( .D(n2500), .CK(clk), .RN(n4375), .Q(
        \key_mem[5][5] ) );
  DFFRX1 \key_mem_reg[9][5]  ( .D(n3012), .CK(clk), .RN(n4431), .Q(
        \key_mem[9][5] ) );
  DFFRX1 \key_mem_reg[5][4]  ( .D(n2501), .CK(clk), .RN(n4412), .Q(
        \key_mem[5][4] ) );
  DFFRX1 \key_mem_reg[9][4]  ( .D(n3013), .CK(clk), .RN(n4467), .Q(
        \key_mem[9][4] ) );
  DFFRX1 \key_mem_reg[5][3]  ( .D(n2502), .CK(clk), .RN(n4381), .Q(
        \key_mem[5][3] ) );
  DFFRX1 \key_mem_reg[9][3]  ( .D(n3014), .CK(clk), .RN(n4385), .Q(
        \key_mem[9][3] ) );
  DFFRX1 \key_mem_reg[5][2]  ( .D(n2503), .CK(clk), .RN(n4374), .Q(
        \key_mem[5][2] ) );
  DFFRX1 \key_mem_reg[9][2]  ( .D(n3015), .CK(clk), .RN(n4563), .Q(
        \key_mem[9][2] ) );
  DFFRX1 \key_mem_reg[5][1]  ( .D(n2504), .CK(clk), .RN(n4564), .Q(
        \key_mem[5][1] ) );
  DFFRX1 \key_mem_reg[9][1]  ( .D(n3016), .CK(clk), .RN(n4554), .Q(
        \key_mem[9][1] ) );
  DFFRX1 \key_mem_reg[5][0]  ( .D(n2505), .CK(clk), .RN(n4556), .Q(
        \key_mem[5][0] ) );
  DFFRX1 \key_mem_reg[9][0]  ( .D(n3017), .CK(clk), .RN(n4556), .Q(
        \key_mem[9][0] ) );
  DFFRX1 \key_mem_reg[5][127]  ( .D(n2378), .CK(clk), .RN(n4527), .Q(
        \key_mem[5][127] ) );
  DFFRX1 \key_mem_reg[9][127]  ( .D(n2890), .CK(clk), .RN(n4534), .Q(
        \key_mem[9][127] ) );
  DFFRX1 \key_mem_reg[5][95]  ( .D(n2410), .CK(clk), .RN(n4563), .Q(
        \key_mem[5][95] ) );
  DFFRX1 \key_mem_reg[9][95]  ( .D(n2922), .CK(clk), .RN(n4515), .Q(
        \key_mem[9][95] ) );
  DFFRX1 \key_mem_reg[5][63]  ( .D(n2442), .CK(clk), .RN(n4505), .Q(
        \key_mem[5][63] ) );
  DFFRX1 \key_mem_reg[9][63]  ( .D(n2954), .CK(clk), .RN(n4514), .Q(
        \key_mem[9][63] ) );
  DFFRX1 \key_mem_reg[5][31]  ( .D(n2474), .CK(clk), .RN(n4557), .Q(
        \key_mem[5][31] ) );
  DFFRX1 \key_mem_reg[9][31]  ( .D(n2986), .CK(clk), .RN(n4557), .Q(
        \key_mem[9][31] ) );
  DFFRX1 \key_mem_reg[5][120]  ( .D(n2385), .CK(clk), .RN(n4493), .Q(
        \key_mem[5][120] ) );
  DFFRX1 \key_mem_reg[9][120]  ( .D(n2897), .CK(clk), .RN(n4492), .Q(
        \key_mem[9][120] ) );
  DFFRX1 \key_mem_reg[5][88]  ( .D(n2417), .CK(clk), .RN(n4558), .Q(
        \key_mem[5][88] ) );
  DFFRX1 \key_mem_reg[9][88]  ( .D(n2929), .CK(clk), .RN(n4558), .Q(
        \key_mem[9][88] ) );
  DFFRX1 \key_mem_reg[5][56]  ( .D(n2449), .CK(clk), .RN(n4476), .Q(
        \key_mem[5][56] ) );
  DFFRX1 \key_mem_reg[9][56]  ( .D(n2961), .CK(clk), .RN(n4512), .Q(
        \key_mem[9][56] ) );
  DFFRX1 \key_mem_reg[5][24]  ( .D(n2481), .CK(clk), .RN(n4454), .Q(
        \key_mem[5][24] ) );
  DFFRX1 \key_mem_reg[9][24]  ( .D(n2993), .CK(clk), .RN(n4554), .Q(
        \key_mem[9][24] ) );
  DFFRX1 \key_mem_reg[5][122]  ( .D(n2383), .CK(clk), .RN(n4485), .Q(
        \key_mem[5][122] ) );
  DFFRX1 \key_mem_reg[9][122]  ( .D(n2895), .CK(clk), .RN(n4486), .Q(
        \key_mem[9][122] ) );
  DFFRX1 \key_mem_reg[5][90]  ( .D(n2415), .CK(clk), .RN(n4487), .Q(
        \key_mem[5][90] ) );
  DFFRX1 \key_mem_reg[9][90]  ( .D(n2927), .CK(clk), .RN(n4487), .Q(
        \key_mem[9][90] ) );
  DFFRX1 \key_mem_reg[5][58]  ( .D(n2447), .CK(clk), .RN(n4489), .Q(
        \key_mem[5][58] ) );
  DFFRX1 \key_mem_reg[9][58]  ( .D(n2959), .CK(clk), .RN(n4489), .Q(
        \key_mem[9][58] ) );
  DFFRX1 \key_mem_reg[5][26]  ( .D(n2479), .CK(clk), .RN(n4490), .Q(
        \key_mem[5][26] ) );
  DFFRX1 \key_mem_reg[9][26]  ( .D(n2991), .CK(clk), .RN(n4491), .Q(
        \key_mem[9][26] ) );
  DFFRX1 \key_mem_reg[5][123]  ( .D(n2382), .CK(clk), .RN(n4484), .Q(
        \key_mem[5][123] ) );
  DFFRX1 \key_mem_reg[9][123]  ( .D(n2894), .CK(clk), .RN(n4433), .Q(
        \key_mem[9][123] ) );
  DFFRX1 \key_mem_reg[5][91]  ( .D(n2414), .CK(clk), .RN(n4492), .Q(
        \key_mem[5][91] ) );
  DFFRX1 \key_mem_reg[9][91]  ( .D(n2926), .CK(clk), .RN(n4493), .Q(
        \key_mem[9][91] ) );
  DFFRX1 \key_mem_reg[5][59]  ( .D(n2446), .CK(clk), .RN(n4494), .Q(
        \key_mem[5][59] ) );
  DFFRX1 \key_mem_reg[9][59]  ( .D(n2958), .CK(clk), .RN(n4494), .Q(
        \key_mem[9][59] ) );
  DFFRX1 \key_mem_reg[5][27]  ( .D(n2478), .CK(clk), .RN(n4496), .Q(
        \key_mem[5][27] ) );
  DFFRX1 \key_mem_reg[9][27]  ( .D(n2990), .CK(clk), .RN(n4470), .Q(
        \key_mem[9][27] ) );
  DFFRX1 \key_mem_reg[5][126]  ( .D(n2379), .CK(clk), .RN(n4471), .Q(
        \key_mem[5][126] ) );
  DFFRX1 \key_mem_reg[9][126]  ( .D(n2891), .CK(clk), .RN(n4472), .Q(
        \key_mem[9][126] ) );
  DFFRX1 \key_mem_reg[5][94]  ( .D(n2411), .CK(clk), .RN(n4473), .Q(
        \key_mem[5][94] ) );
  DFFRX1 \key_mem_reg[9][94]  ( .D(n2923), .CK(clk), .RN(n4474), .Q(
        \key_mem[9][94] ) );
  DFFRX1 \key_mem_reg[5][62]  ( .D(n2443), .CK(clk), .RN(n4475), .Q(
        \key_mem[5][62] ) );
  DFFRX1 \key_mem_reg[9][62]  ( .D(n2955), .CK(clk), .RN(n4475), .Q(
        \key_mem[9][62] ) );
  DFFRX1 \key_mem_reg[5][30]  ( .D(n2475), .CK(clk), .RN(n4477), .Q(
        \key_mem[5][30] ) );
  DFFRX1 \key_mem_reg[9][30]  ( .D(n2987), .CK(clk), .RN(n4477), .Q(
        \key_mem[9][30] ) );
  DFFRX1 \key_mem_reg[5][125]  ( .D(n2380), .CK(clk), .RN(n4479), .Q(
        \key_mem[5][125] ) );
  DFFRX1 \key_mem_reg[9][125]  ( .D(n2892), .CK(clk), .RN(n4479), .Q(
        \key_mem[9][125] ) );
  DFFRX1 \key_mem_reg[5][93]  ( .D(n2412), .CK(clk), .RN(n4480), .Q(
        \key_mem[5][93] ) );
  DFFRX1 \key_mem_reg[9][93]  ( .D(n2924), .CK(clk), .RN(n4481), .Q(
        \key_mem[9][93] ) );
  DFFRX1 \key_mem_reg[5][61]  ( .D(n2444), .CK(clk), .RN(n4482), .Q(
        \key_mem[5][61] ) );
  DFFRX1 \key_mem_reg[9][61]  ( .D(n2956), .CK(clk), .RN(n4483), .Q(
        \key_mem[9][61] ) );
  DFFRX1 \key_mem_reg[5][29]  ( .D(n2476), .CK(clk), .RN(n4484), .Q(
        \key_mem[5][29] ) );
  DFFRX1 \key_mem_reg[9][29]  ( .D(n2988), .CK(clk), .RN(n4484), .Q(
        \key_mem[9][29] ) );
  DFFRX1 \key_mem_reg[5][124]  ( .D(n2381), .CK(clk), .RN(n4512), .Q(
        \key_mem[5][124] ) );
  DFFRX1 \key_mem_reg[9][124]  ( .D(n2893), .CK(clk), .RN(n4512), .Q(
        \key_mem[9][124] ) );
  DFFRX1 \key_mem_reg[5][92]  ( .D(n2413), .CK(clk), .RN(n4513), .Q(
        \key_mem[5][92] ) );
  DFFRX1 \key_mem_reg[9][92]  ( .D(n2925), .CK(clk), .RN(n4514), .Q(
        \key_mem[9][92] ) );
  DFFRX1 \key_mem_reg[5][60]  ( .D(n2445), .CK(clk), .RN(n4515), .Q(
        \key_mem[5][60] ) );
  DFFRX1 \key_mem_reg[9][60]  ( .D(n2957), .CK(clk), .RN(n4516), .Q(
        \key_mem[9][60] ) );
  DFFRX1 \key_mem_reg[5][28]  ( .D(n2477), .CK(clk), .RN(n4517), .Q(
        \key_mem[5][28] ) );
  DFFRX1 \key_mem_reg[9][28]  ( .D(n2989), .CK(clk), .RN(n4517), .Q(
        \key_mem[9][28] ) );
  DFFRX1 \key_mem_reg[5][121]  ( .D(n2384), .CK(clk), .RN(n4519), .Q(
        \key_mem[5][121] ) );
  DFFRX1 \key_mem_reg[9][121]  ( .D(n2896), .CK(clk), .RN(n4519), .Q(
        \key_mem[9][121] ) );
  DFFRX1 \key_mem_reg[5][89]  ( .D(n2416), .CK(clk), .RN(n4521), .Q(
        \key_mem[5][89] ) );
  DFFRX1 \key_mem_reg[9][89]  ( .D(n2928), .CK(clk), .RN(n4521), .Q(
        \key_mem[9][89] ) );
  DFFRX1 \key_mem_reg[5][57]  ( .D(n2448), .CK(clk), .RN(n4522), .Q(
        \key_mem[5][57] ) );
  DFFRX1 \key_mem_reg[9][57]  ( .D(n2960), .CK(clk), .RN(n4523), .Q(
        \key_mem[9][57] ) );
  DFFRX1 \key_mem_reg[5][25]  ( .D(n2480), .CK(clk), .RN(n4524), .Q(
        \key_mem[5][25] ) );
  DFFRX1 \key_mem_reg[9][25]  ( .D(n2992), .CK(clk), .RN(n4525), .Q(
        \key_mem[9][25] ) );
  DFFRX1 \key_mem_reg[1][127]  ( .D(n1866), .CK(clk), .RN(n4525), .Q(
        \key_mem[1][127] ) );
  DFFRX1 \key_mem_reg[1][126]  ( .D(n1867), .CK(clk), .RN(n4525), .Q(
        \key_mem[1][126] ) );
  DFFRX1 \key_mem_reg[1][125]  ( .D(n1868), .CK(clk), .RN(n4526), .Q(
        \key_mem[1][125] ) );
  DFFRX1 \key_mem_reg[1][124]  ( .D(n1869), .CK(clk), .RN(n4526), .Q(
        \key_mem[1][124] ) );
  DFFRX1 \key_mem_reg[1][123]  ( .D(n1870), .CK(clk), .RN(n4526), .Q(
        \key_mem[1][123] ) );
  DFFRX1 \key_mem_reg[1][122]  ( .D(n1871), .CK(clk), .RN(n4526), .Q(
        \key_mem[1][122] ) );
  DFFRX1 \key_mem_reg[1][121]  ( .D(n1872), .CK(clk), .RN(n4503), .Q(
        \key_mem[1][121] ) );
  DFFRX1 \key_mem_reg[1][120]  ( .D(n1873), .CK(clk), .RN(n4496), .Q(
        \key_mem[1][120] ) );
  DFFRX1 \key_mem_reg[1][119]  ( .D(n1874), .CK(clk), .RN(n4496), .Q(
        \key_mem[1][119] ) );
  DFFRX1 \key_mem_reg[1][118]  ( .D(n1875), .CK(clk), .RN(n4496), .Q(
        \key_mem[1][118] ) );
  DFFRX1 \key_mem_reg[1][117]  ( .D(n1876), .CK(clk), .RN(n4496), .Q(
        \key_mem[1][117] ) );
  DFFRX1 \key_mem_reg[1][116]  ( .D(n1877), .CK(clk), .RN(n4496), .Q(
        \key_mem[1][116] ) );
  DFFRX1 \key_mem_reg[1][115]  ( .D(n1878), .CK(clk), .RN(n4497), .Q(
        \key_mem[1][115] ) );
  DFFRX1 \key_mem_reg[1][114]  ( .D(n1879), .CK(clk), .RN(n4497), .Q(
        \key_mem[1][114] ) );
  DFFRX1 \key_mem_reg[1][113]  ( .D(n1880), .CK(clk), .RN(n4497), .Q(
        \key_mem[1][113] ) );
  DFFRX1 \key_mem_reg[1][112]  ( .D(n1881), .CK(clk), .RN(n4497), .Q(
        \key_mem[1][112] ) );
  DFFRX1 \key_mem_reg[1][111]  ( .D(n1882), .CK(clk), .RN(n4497), .Q(
        \key_mem[1][111] ) );
  DFFRX1 \key_mem_reg[1][110]  ( .D(n1883), .CK(clk), .RN(n4497), .Q(
        \key_mem[1][110] ) );
  DFFRX1 \key_mem_reg[1][109]  ( .D(n1884), .CK(clk), .RN(n4497), .Q(
        \key_mem[1][109] ) );
  DFFRX1 \key_mem_reg[1][108]  ( .D(n1885), .CK(clk), .RN(n4497), .Q(
        \key_mem[1][108] ) );
  DFFRX1 \key_mem_reg[1][107]  ( .D(n1886), .CK(clk), .RN(n4498), .Q(
        \key_mem[1][107] ) );
  DFFRX1 \key_mem_reg[1][106]  ( .D(n1887), .CK(clk), .RN(n4498), .Q(
        \key_mem[1][106] ) );
  DFFRX1 \key_mem_reg[1][105]  ( .D(n1888), .CK(clk), .RN(n4498), .Q(
        \key_mem[1][105] ) );
  DFFRX1 \key_mem_reg[1][104]  ( .D(n1889), .CK(clk), .RN(n4498), .Q(
        \key_mem[1][104] ) );
  DFFRX1 \key_mem_reg[1][103]  ( .D(n1890), .CK(clk), .RN(n4498), .Q(
        \key_mem[1][103] ) );
  DFFRX1 \key_mem_reg[1][102]  ( .D(n1891), .CK(clk), .RN(n4498), .Q(
        \key_mem[1][102] ) );
  DFFRX1 \key_mem_reg[1][101]  ( .D(n1892), .CK(clk), .RN(n4498), .Q(
        \key_mem[1][101] ) );
  DFFRX1 \key_mem_reg[1][100]  ( .D(n1893), .CK(clk), .RN(n4498), .Q(
        \key_mem[1][100] ) );
  DFFRX1 \key_mem_reg[1][99]  ( .D(n1894), .CK(clk), .RN(n4499), .Q(
        \key_mem[1][99] ) );
  DFFRX1 \key_mem_reg[1][98]  ( .D(n1895), .CK(clk), .RN(n4499), .Q(
        \key_mem[1][98] ) );
  DFFRX1 \key_mem_reg[1][97]  ( .D(n1896), .CK(clk), .RN(n4499), .Q(
        \key_mem[1][97] ) );
  DFFRX1 \key_mem_reg[1][96]  ( .D(n1897), .CK(clk), .RN(n4499), .Q(
        \key_mem[1][96] ) );
  DFFRX1 \key_mem_reg[1][95]  ( .D(n1898), .CK(clk), .RN(n4499), .Q(
        \key_mem[1][95] ) );
  DFFRX1 \key_mem_reg[1][94]  ( .D(n1899), .CK(clk), .RN(n4499), .Q(
        \key_mem[1][94] ) );
  DFFRX1 \key_mem_reg[1][93]  ( .D(n1900), .CK(clk), .RN(n4499), .Q(
        \key_mem[1][93] ) );
  DFFRX1 \key_mem_reg[1][92]  ( .D(n1901), .CK(clk), .RN(n4499), .Q(
        \key_mem[1][92] ) );
  DFFRX1 \key_mem_reg[1][91]  ( .D(n1902), .CK(clk), .RN(n4500), .Q(
        \key_mem[1][91] ) );
  DFFRX1 \key_mem_reg[1][90]  ( .D(n1903), .CK(clk), .RN(n4500), .Q(
        \key_mem[1][90] ) );
  DFFRX1 \key_mem_reg[1][89]  ( .D(n1904), .CK(clk), .RN(n4500), .Q(
        \key_mem[1][89] ) );
  DFFRX1 \key_mem_reg[1][88]  ( .D(n1905), .CK(clk), .RN(n4500), .Q(
        \key_mem[1][88] ) );
  DFFRX1 \key_mem_reg[1][87]  ( .D(n1906), .CK(clk), .RN(n4500), .Q(
        \key_mem[1][87] ) );
  DFFRX1 \key_mem_reg[1][86]  ( .D(n1907), .CK(clk), .RN(n4500), .Q(
        \key_mem[1][86] ) );
  DFFRX1 \key_mem_reg[1][85]  ( .D(n1908), .CK(clk), .RN(n4500), .Q(
        \key_mem[1][85] ) );
  DFFRX1 \key_mem_reg[1][84]  ( .D(n1909), .CK(clk), .RN(n4500), .Q(
        \key_mem[1][84] ) );
  DFFRX1 \key_mem_reg[1][83]  ( .D(n1910), .CK(clk), .RN(n4501), .Q(
        \key_mem[1][83] ) );
  DFFRX1 \key_mem_reg[1][82]  ( .D(n1911), .CK(clk), .RN(n4501), .Q(
        \key_mem[1][82] ) );
  DFFRX1 \key_mem_reg[1][81]  ( .D(n1912), .CK(clk), .RN(n4501), .Q(
        \key_mem[1][81] ) );
  DFFRX1 \key_mem_reg[1][80]  ( .D(n1913), .CK(clk), .RN(n4501), .Q(
        \key_mem[1][80] ) );
  DFFRX1 \key_mem_reg[1][79]  ( .D(n1914), .CK(clk), .RN(n4501), .Q(
        \key_mem[1][79] ) );
  DFFRX1 \key_mem_reg[1][78]  ( .D(n1915), .CK(clk), .RN(n4501), .Q(
        \key_mem[1][78] ) );
  DFFRX1 \key_mem_reg[1][77]  ( .D(n1916), .CK(clk), .RN(n4501), .Q(
        \key_mem[1][77] ) );
  DFFRX1 \key_mem_reg[1][76]  ( .D(n1917), .CK(clk), .RN(n4501), .Q(
        \key_mem[1][76] ) );
  DFFRX1 \key_mem_reg[1][75]  ( .D(n1918), .CK(clk), .RN(n4502), .Q(
        \key_mem[1][75] ) );
  DFFRX1 \key_mem_reg[1][74]  ( .D(n1919), .CK(clk), .RN(n4502), .Q(
        \key_mem[1][74] ) );
  DFFRX1 \key_mem_reg[1][73]  ( .D(n1920), .CK(clk), .RN(n4502), .Q(
        \key_mem[1][73] ) );
  DFFRX1 \key_mem_reg[1][72]  ( .D(n1921), .CK(clk), .RN(n4502), .Q(
        \key_mem[1][72] ) );
  DFFRX1 \key_mem_reg[1][71]  ( .D(n1922), .CK(clk), .RN(n4502), .Q(
        \key_mem[1][71] ) );
  DFFRX1 \key_mem_reg[1][70]  ( .D(n1923), .CK(clk), .RN(n4502), .Q(
        \key_mem[1][70] ) );
  DFFRX1 \key_mem_reg[1][69]  ( .D(n1924), .CK(clk), .RN(n4502), .Q(
        \key_mem[1][69] ) );
  DFFRX1 \key_mem_reg[1][68]  ( .D(n1925), .CK(clk), .RN(n4502), .Q(
        \key_mem[1][68] ) );
  DFFRX1 \key_mem_reg[1][67]  ( .D(n1926), .CK(clk), .RN(n4503), .Q(
        \key_mem[1][67] ) );
  DFFRX1 \key_mem_reg[1][66]  ( .D(n1927), .CK(clk), .RN(n4503), .Q(
        \key_mem[1][66] ) );
  DFFRX1 \key_mem_reg[1][65]  ( .D(n1928), .CK(clk), .RN(n4503), .Q(
        \key_mem[1][65] ) );
  DFFRX1 \key_mem_reg[1][64]  ( .D(n1929), .CK(clk), .RN(n4503), .Q(
        \key_mem[1][64] ) );
  DFFRX1 \key_mem_reg[1][63]  ( .D(n1930), .CK(clk), .RN(n4503), .Q(
        \key_mem[1][63] ) );
  DFFRX1 \key_mem_reg[1][62]  ( .D(n1931), .CK(clk), .RN(n4503), .Q(
        \key_mem[1][62] ) );
  DFFRX1 \key_mem_reg[1][61]  ( .D(n1932), .CK(clk), .RN(n4503), .Q(
        \key_mem[1][61] ) );
  DFFRX1 \key_mem_reg[1][60]  ( .D(n1933), .CK(clk), .RN(n4504), .Q(
        \key_mem[1][60] ) );
  DFFRX1 \key_mem_reg[1][59]  ( .D(n1934), .CK(clk), .RN(n4504), .Q(
        \key_mem[1][59] ) );
  DFFRX1 \key_mem_reg[1][58]  ( .D(n1935), .CK(clk), .RN(n4504), .Q(
        \key_mem[1][58] ) );
  DFFRX1 \key_mem_reg[1][57]  ( .D(n1936), .CK(clk), .RN(n4504), .Q(
        \key_mem[1][57] ) );
  DFFRX1 \key_mem_reg[1][56]  ( .D(n1937), .CK(clk), .RN(n4504), .Q(
        \key_mem[1][56] ) );
  DFFRX1 \key_mem_reg[1][55]  ( .D(n1938), .CK(clk), .RN(n4504), .Q(
        \key_mem[1][55] ) );
  DFFRX1 \key_mem_reg[1][54]  ( .D(n1939), .CK(clk), .RN(n4504), .Q(
        \key_mem[1][54] ) );
  DFFRX1 \key_mem_reg[1][53]  ( .D(n1940), .CK(clk), .RN(n4504), .Q(
        \key_mem[1][53] ) );
  DFFRX1 \key_mem_reg[1][52]  ( .D(n1941), .CK(clk), .RN(n4505), .Q(
        \key_mem[1][52] ) );
  DFFRX1 \key_mem_reg[1][51]  ( .D(n1942), .CK(clk), .RN(n4505), .Q(
        \key_mem[1][51] ) );
  DFFRX1 \key_mem_reg[1][50]  ( .D(n1943), .CK(clk), .RN(n4505), .Q(
        \key_mem[1][50] ) );
  DFFRX1 \key_mem_reg[1][49]  ( .D(n1944), .CK(clk), .RN(n4505), .Q(
        \key_mem[1][49] ) );
  DFFRX1 \key_mem_reg[1][47]  ( .D(n1946), .CK(clk), .RN(n4505), .Q(
        \key_mem[1][47] ) );
  DFFRX1 \key_mem_reg[1][46]  ( .D(n1947), .CK(clk), .RN(n4505), .Q(
        \key_mem[1][46] ) );
  DFFRX1 \key_mem_reg[1][45]  ( .D(n1948), .CK(clk), .RN(n4505), .Q(
        \key_mem[1][45] ) );
  DFFRX1 \key_mem_reg[1][44]  ( .D(n1949), .CK(clk), .RN(n4506), .Q(
        \key_mem[1][44] ) );
  DFFRX1 \key_mem_reg[1][43]  ( .D(n1950), .CK(clk), .RN(n4506), .Q(
        \key_mem[1][43] ) );
  DFFRX1 \key_mem_reg[1][42]  ( .D(n1951), .CK(clk), .RN(n4506), .Q(
        \key_mem[1][42] ) );
  DFFRX1 \key_mem_reg[1][41]  ( .D(n1952), .CK(clk), .RN(n4506), .Q(
        \key_mem[1][41] ) );
  DFFRX1 \key_mem_reg[1][40]  ( .D(n1953), .CK(clk), .RN(n4506), .Q(
        \key_mem[1][40] ) );
  DFFRX1 \key_mem_reg[1][39]  ( .D(n1954), .CK(clk), .RN(n4506), .Q(
        \key_mem[1][39] ) );
  DFFRX1 \key_mem_reg[1][38]  ( .D(n1955), .CK(clk), .RN(n4506), .Q(
        \key_mem[1][38] ) );
  DFFRX1 \key_mem_reg[1][37]  ( .D(n1956), .CK(clk), .RN(n4506), .Q(
        \key_mem[1][37] ) );
  DFFRX1 \key_mem_reg[1][36]  ( .D(n1957), .CK(clk), .RN(n4507), .Q(
        \key_mem[1][36] ) );
  DFFRX1 \key_mem_reg[1][35]  ( .D(n1958), .CK(clk), .RN(n4507), .Q(
        \key_mem[1][35] ) );
  DFFRX1 \key_mem_reg[1][34]  ( .D(n1959), .CK(clk), .RN(n4507), .Q(
        \key_mem[1][34] ) );
  DFFRX1 \key_mem_reg[1][33]  ( .D(n1960), .CK(clk), .RN(n4507), .Q(
        \key_mem[1][33] ) );
  DFFRX1 \key_mem_reg[1][32]  ( .D(n1961), .CK(clk), .RN(n4507), .Q(
        \key_mem[1][32] ) );
  DFFRX1 \key_mem_reg[1][31]  ( .D(n1962), .CK(clk), .RN(n4507), .Q(
        \key_mem[1][31] ) );
  DFFRX1 \key_mem_reg[1][30]  ( .D(n1963), .CK(clk), .RN(n4507), .Q(
        \key_mem[1][30] ) );
  DFFRX1 \key_mem_reg[1][29]  ( .D(n1964), .CK(clk), .RN(n4507), .Q(
        \key_mem[1][29] ) );
  DFFRX1 \key_mem_reg[1][28]  ( .D(n1965), .CK(clk), .RN(n4508), .Q(
        \key_mem[1][28] ) );
  DFFRX1 \key_mem_reg[1][27]  ( .D(n1966), .CK(clk), .RN(n4508), .Q(
        \key_mem[1][27] ) );
  DFFRX1 \key_mem_reg[1][26]  ( .D(n1967), .CK(clk), .RN(n4508), .Q(
        \key_mem[1][26] ) );
  DFFRX1 \key_mem_reg[1][25]  ( .D(n1968), .CK(clk), .RN(n4508), .Q(
        \key_mem[1][25] ) );
  DFFRX1 \key_mem_reg[1][24]  ( .D(n1969), .CK(clk), .RN(n4508), .Q(
        \key_mem[1][24] ) );
  DFFRX1 \key_mem_reg[1][23]  ( .D(n1970), .CK(clk), .RN(n4508), .Q(
        \key_mem[1][23] ) );
  DFFRX1 \key_mem_reg[1][22]  ( .D(n1971), .CK(clk), .RN(n4508), .Q(
        \key_mem[1][22] ) );
  DFFRX1 \key_mem_reg[1][21]  ( .D(n1972), .CK(clk), .RN(n4508), .Q(
        \key_mem[1][21] ) );
  DFFRX1 \key_mem_reg[1][20]  ( .D(n1973), .CK(clk), .RN(n4509), .Q(
        \key_mem[1][20] ) );
  DFFRX1 \key_mem_reg[1][19]  ( .D(n1974), .CK(clk), .RN(n4509), .Q(
        \key_mem[1][19] ) );
  DFFRX1 \key_mem_reg[1][18]  ( .D(n1975), .CK(clk), .RN(n4509), .Q(
        \key_mem[1][18] ) );
  DFFRX1 \key_mem_reg[1][17]  ( .D(n1976), .CK(clk), .RN(n4509), .Q(
        \key_mem[1][17] ) );
  DFFRX1 \key_mem_reg[1][16]  ( .D(n1977), .CK(clk), .RN(n4509), .Q(
        \key_mem[1][16] ) );
  DFFRX1 \key_mem_reg[1][15]  ( .D(n1978), .CK(clk), .RN(n4509), .Q(
        \key_mem[1][15] ) );
  DFFRX1 \key_mem_reg[1][14]  ( .D(n1979), .CK(clk), .RN(n4509), .Q(
        \key_mem[1][14] ) );
  DFFRX1 \key_mem_reg[1][13]  ( .D(n1980), .CK(clk), .RN(n4509), .Q(
        \key_mem[1][13] ) );
  DFFRX1 \key_mem_reg[1][12]  ( .D(n1981), .CK(clk), .RN(n4510), .Q(
        \key_mem[1][12] ) );
  DFFRX1 \key_mem_reg[1][11]  ( .D(n1982), .CK(clk), .RN(n4510), .Q(
        \key_mem[1][11] ) );
  DFFRX1 \key_mem_reg[1][10]  ( .D(n1983), .CK(clk), .RN(n4510), .Q(
        \key_mem[1][10] ) );
  DFFRX1 \key_mem_reg[1][9]  ( .D(n1984), .CK(clk), .RN(n4510), .Q(
        \key_mem[1][9] ) );
  DFFRX1 \key_mem_reg[1][8]  ( .D(n1985), .CK(clk), .RN(n4510), .Q(
        \key_mem[1][8] ) );
  DFFRX1 \key_mem_reg[1][7]  ( .D(n1986), .CK(clk), .RN(n4510), .Q(
        \key_mem[1][7] ) );
  DFFRX1 \key_mem_reg[1][6]  ( .D(n1987), .CK(clk), .RN(n4510), .Q(
        \key_mem[1][6] ) );
  DFFRX1 \key_mem_reg[1][5]  ( .D(n1988), .CK(clk), .RN(n4510), .Q(
        \key_mem[1][5] ) );
  DFFRX1 \key_mem_reg[1][4]  ( .D(n1989), .CK(clk), .RN(n4511), .Q(
        \key_mem[1][4] ) );
  DFFRX1 \key_mem_reg[1][3]  ( .D(n1990), .CK(clk), .RN(n4511), .Q(
        \key_mem[1][3] ) );
  DFFRX1 \key_mem_reg[1][2]  ( .D(n1991), .CK(clk), .RN(n4511), .Q(
        \key_mem[1][2] ) );
  DFFRX1 \key_mem_reg[1][1]  ( .D(n1992), .CK(clk), .RN(n4511), .Q(
        \key_mem[1][1] ) );
  DFFRX1 \key_mem_reg[1][0]  ( .D(n1993), .CK(clk), .RN(n4526), .Q(
        \key_mem[1][0] ) );
  DFFRX1 \key_mem_reg[3][119]  ( .D(n2130), .CK(clk), .RN(n4430), .Q(
        \key_mem[3][119] ) );
  DFFRX1 \key_mem_reg[7][119]  ( .D(n2642), .CK(clk), .RN(n4430), .Q(
        \key_mem[7][119] ) );
  DFFRX1 \key_mem_reg[11][119]  ( .D(n3154), .CK(clk), .RN(n4431), .Q(
        \key_mem[11][119] ) );
  DFFRX1 \key_mem_reg[3][118]  ( .D(n2131), .CK(clk), .RN(n4432), .Q(
        \key_mem[3][118] ) );
  DFFRX1 \key_mem_reg[7][118]  ( .D(n2643), .CK(clk), .RN(n4432), .Q(
        \key_mem[7][118] ) );
  DFFRX1 \key_mem_reg[11][118]  ( .D(n3155), .CK(clk), .RN(n4373), .Q(
        \key_mem[11][118] ) );
  DFFRX1 \key_mem_reg[3][117]  ( .D(n2132), .CK(clk), .RN(n4372), .Q(
        \key_mem[3][117] ) );
  DFFRX1 \key_mem_reg[7][117]  ( .D(n2644), .CK(clk), .RN(n4433), .Q(
        \key_mem[7][117] ) );
  DFFRX1 \key_mem_reg[11][117]  ( .D(n3156), .CK(clk), .RN(n4433), .Q(
        \key_mem[11][117] ) );
  DFFRX1 \key_mem_reg[3][116]  ( .D(n2133), .CK(clk), .RN(n4498), .Q(
        \key_mem[3][116] ) );
  DFFRX1 \key_mem_reg[7][116]  ( .D(n2645), .CK(clk), .RN(n4404), .Q(
        \key_mem[7][116] ) );
  DFFRX1 \key_mem_reg[11][116]  ( .D(n3157), .CK(clk), .RN(n4403), .Q(
        \key_mem[11][116] ) );
  DFFRX1 \key_mem_reg[3][115]  ( .D(n2134), .CK(clk), .RN(n4396), .Q(
        \key_mem[3][115] ) );
  DFFRX1 \key_mem_reg[7][115]  ( .D(n2646), .CK(clk), .RN(n4434), .Q(
        \key_mem[7][115] ) );
  DFFRX1 \key_mem_reg[11][115]  ( .D(n3158), .CK(clk), .RN(n4434), .Q(
        \key_mem[11][115] ) );
  DFFRX1 \key_mem_reg[3][114]  ( .D(n2135), .CK(clk), .RN(n4435), .Q(
        \key_mem[3][114] ) );
  DFFRX1 \key_mem_reg[7][114]  ( .D(n2647), .CK(clk), .RN(n4435), .Q(
        \key_mem[7][114] ) );
  DFFRX1 \key_mem_reg[11][114]  ( .D(n3159), .CK(clk), .RN(n4436), .Q(
        \key_mem[11][114] ) );
  DFFRX1 \key_mem_reg[3][113]  ( .D(n2136), .CK(clk), .RN(n4437), .Q(
        \key_mem[3][113] ) );
  DFFRX1 \key_mem_reg[7][113]  ( .D(n2648), .CK(clk), .RN(n4437), .Q(
        \key_mem[7][113] ) );
  DFFRX1 \key_mem_reg[11][113]  ( .D(n3160), .CK(clk), .RN(n4438), .Q(
        \key_mem[11][113] ) );
  DFFRX1 \key_mem_reg[3][112]  ( .D(n2137), .CK(clk), .RN(n4438), .Q(
        \key_mem[3][112] ) );
  DFFRX1 \key_mem_reg[7][112]  ( .D(n2649), .CK(clk), .RN(n4439), .Q(
        \key_mem[7][112] ) );
  DFFRX1 \key_mem_reg[11][112]  ( .D(n3161), .CK(clk), .RN(n4439), .Q(
        \key_mem[11][112] ) );
  DFFRX1 \key_mem_reg[3][111]  ( .D(n2138), .CK(clk), .RN(n4440), .Q(
        \key_mem[3][111] ) );
  DFFRX1 \key_mem_reg[7][111]  ( .D(n2650), .CK(clk), .RN(n4417), .Q(
        \key_mem[7][111] ) );
  DFFRX1 \key_mem_reg[11][111]  ( .D(n3162), .CK(clk), .RN(n4418), .Q(
        \key_mem[11][111] ) );
  DFFRX1 \key_mem_reg[3][110]  ( .D(n2139), .CK(clk), .RN(n4440), .Q(
        \key_mem[3][110] ) );
  DFFRX1 \key_mem_reg[7][110]  ( .D(n2651), .CK(clk), .RN(n4437), .Q(
        \key_mem[7][110] ) );
  DFFRX1 \key_mem_reg[11][110]  ( .D(n3163), .CK(clk), .RN(n4419), .Q(
        \key_mem[11][110] ) );
  DFFRX1 \key_mem_reg[3][109]  ( .D(n2140), .CK(clk), .RN(n4419), .Q(
        \key_mem[3][109] ) );
  DFFRX1 \key_mem_reg[7][109]  ( .D(n2652), .CK(clk), .RN(n4420), .Q(
        \key_mem[7][109] ) );
  DFFRX1 \key_mem_reg[11][109]  ( .D(n3164), .CK(clk), .RN(n4420), .Q(
        \key_mem[11][109] ) );
  DFFRX1 \key_mem_reg[3][108]  ( .D(n2141), .CK(clk), .RN(n4421), .Q(
        \key_mem[3][108] ) );
  DFFRX1 \key_mem_reg[7][108]  ( .D(n2653), .CK(clk), .RN(n4422), .Q(
        \key_mem[7][108] ) );
  DFFRX1 \key_mem_reg[11][108]  ( .D(n3165), .CK(clk), .RN(n4422), .Q(
        \key_mem[11][108] ) );
  DFFRX1 \key_mem_reg[3][106]  ( .D(n2143), .CK(clk), .RN(n4423), .Q(
        \key_mem[3][106] ) );
  DFFRX1 \key_mem_reg[7][106]  ( .D(n2655), .CK(clk), .RN(n4423), .Q(
        \key_mem[7][106] ) );
  DFFRX1 \key_mem_reg[11][106]  ( .D(n3167), .CK(clk), .RN(n4424), .Q(
        \key_mem[11][106] ) );
  DFFRX1 \key_mem_reg[3][105]  ( .D(n2144), .CK(clk), .RN(n4424), .Q(
        \key_mem[3][105] ) );
  DFFRX1 \key_mem_reg[7][105]  ( .D(n2656), .CK(clk), .RN(n4425), .Q(
        \key_mem[7][105] ) );
  DFFRX1 \key_mem_reg[11][105]  ( .D(n3168), .CK(clk), .RN(n4425), .Q(
        \key_mem[11][105] ) );
  DFFRX1 \key_mem_reg[3][104]  ( .D(n2145), .CK(clk), .RN(n4426), .Q(
        \key_mem[3][104] ) );
  DFFRX1 \key_mem_reg[7][104]  ( .D(n2657), .CK(clk), .RN(n4427), .Q(
        \key_mem[7][104] ) );
  DFFRX1 \key_mem_reg[11][104]  ( .D(n3169), .CK(clk), .RN(n4427), .Q(
        \key_mem[11][104] ) );
  DFFRX1 \key_mem_reg[3][103]  ( .D(n2146), .CK(clk), .RN(n4428), .Q(
        \key_mem[3][103] ) );
  DFFRX1 \key_mem_reg[7][103]  ( .D(n2658), .CK(clk), .RN(n4428), .Q(
        \key_mem[7][103] ) );
  DFFRX1 \key_mem_reg[11][103]  ( .D(n3170), .CK(clk), .RN(n4429), .Q(
        \key_mem[11][103] ) );
  DFFRX1 \key_mem_reg[3][102]  ( .D(n2147), .CK(clk), .RN(n4456), .Q(
        \key_mem[3][102] ) );
  DFFRX1 \key_mem_reg[7][102]  ( .D(n2659), .CK(clk), .RN(n4456), .Q(
        \key_mem[7][102] ) );
  DFFRX1 \key_mem_reg[11][102]  ( .D(n3171), .CK(clk), .RN(n4457), .Q(
        \key_mem[11][102] ) );
  DFFRX1 \key_mem_reg[3][101]  ( .D(n2148), .CK(clk), .RN(n4458), .Q(
        \key_mem[3][101] ) );
  DFFRX1 \key_mem_reg[7][101]  ( .D(n2660), .CK(clk), .RN(n4458), .Q(
        \key_mem[7][101] ) );
  DFFRX1 \key_mem_reg[11][101]  ( .D(n3172), .CK(clk), .RN(n4459), .Q(
        \key_mem[11][101] ) );
  DFFRX1 \key_mem_reg[3][100]  ( .D(n2149), .CK(clk), .RN(n4459), .Q(
        \key_mem[3][100] ) );
  DFFRX1 \key_mem_reg[7][100]  ( .D(n2661), .CK(clk), .RN(n4460), .Q(
        \key_mem[7][100] ) );
  DFFRX1 \key_mem_reg[11][100]  ( .D(n3173), .CK(clk), .RN(n4460), .Q(
        \key_mem[11][100] ) );
  DFFRX1 \key_mem_reg[3][99]  ( .D(n2150), .CK(clk), .RN(n4468), .Q(
        \key_mem[3][99] ) );
  DFFRX1 \key_mem_reg[7][99]  ( .D(n2662), .CK(clk), .RN(n4461), .Q(
        \key_mem[7][99] ) );
  DFFRX1 \key_mem_reg[11][99]  ( .D(n3174), .CK(clk), .RN(n4461), .Q(
        \key_mem[11][99] ) );
  DFFRX1 \key_mem_reg[3][98]  ( .D(n2151), .CK(clk), .RN(n4462), .Q(
        \key_mem[3][98] ) );
  DFFRX1 \key_mem_reg[7][98]  ( .D(n2663), .CK(clk), .RN(n4462), .Q(
        \key_mem[7][98] ) );
  DFFRX1 \key_mem_reg[11][98]  ( .D(n3175), .CK(clk), .RN(n4463), .Q(
        \key_mem[11][98] ) );
  DFFRX1 \key_mem_reg[3][97]  ( .D(n2152), .CK(clk), .RN(n4464), .Q(
        \key_mem[3][97] ) );
  DFFRX1 \key_mem_reg[7][97]  ( .D(n2664), .CK(clk), .RN(n4464), .Q(
        \key_mem[7][97] ) );
  DFFRX1 \key_mem_reg[11][97]  ( .D(n3176), .CK(clk), .RN(n4465), .Q(
        \key_mem[11][97] ) );
  DFFRX1 \key_mem_reg[3][96]  ( .D(n2153), .CK(clk), .RN(n4465), .Q(
        \key_mem[3][96] ) );
  DFFRX1 \key_mem_reg[7][96]  ( .D(n2665), .CK(clk), .RN(n4466), .Q(
        \key_mem[7][96] ) );
  DFFRX1 \key_mem_reg[11][96]  ( .D(n3177), .CK(clk), .RN(n4466), .Q(
        \key_mem[11][96] ) );
  DFFRX1 \key_mem_reg[3][87]  ( .D(n2162), .CK(clk), .RN(n4467), .Q(
        \key_mem[3][87] ) );
  DFFRX1 \key_mem_reg[7][87]  ( .D(n2674), .CK(clk), .RN(n4468), .Q(
        \key_mem[7][87] ) );
  DFFRX1 \key_mem_reg[11][87]  ( .D(n3186), .CK(clk), .RN(n4468), .Q(
        \key_mem[11][87] ) );
  DFFRX1 \key_mem_reg[3][86]  ( .D(n2163), .CK(clk), .RN(n4469), .Q(
        \key_mem[3][86] ) );
  DFFRX1 \key_mem_reg[7][86]  ( .D(n2675), .CK(clk), .RN(n4469), .Q(
        \key_mem[7][86] ) );
  DFFRX1 \key_mem_reg[11][86]  ( .D(n3187), .CK(clk), .RN(n4441), .Q(
        \key_mem[11][86] ) );
  DFFRX1 \key_mem_reg[3][85]  ( .D(n2164), .CK(clk), .RN(n4441), .Q(
        \key_mem[3][85] ) );
  DFFRX1 \key_mem_reg[7][85]  ( .D(n2676), .CK(clk), .RN(n4442), .Q(
        \key_mem[7][85] ) );
  DFFRX1 \key_mem_reg[11][85]  ( .D(n3188), .CK(clk), .RN(n4442), .Q(
        \key_mem[11][85] ) );
  DFFRX1 \key_mem_reg[3][84]  ( .D(n2165), .CK(clk), .RN(n4443), .Q(
        \key_mem[3][84] ) );
  DFFRX1 \key_mem_reg[7][84]  ( .D(n2677), .CK(clk), .RN(n4444), .Q(
        \key_mem[7][84] ) );
  DFFRX1 \key_mem_reg[11][84]  ( .D(n3189), .CK(clk), .RN(n4444), .Q(
        \key_mem[11][84] ) );
  DFFRX1 \key_mem_reg[3][83]  ( .D(n2166), .CK(clk), .RN(n4445), .Q(
        \key_mem[3][83] ) );
  DFFRX1 \key_mem_reg[7][83]  ( .D(n2678), .CK(clk), .RN(n4445), .Q(
        \key_mem[7][83] ) );
  DFFRX1 \key_mem_reg[11][83]  ( .D(n3190), .CK(clk), .RN(n4446), .Q(
        \key_mem[11][83] ) );
  DFFRX1 \key_mem_reg[3][82]  ( .D(n2167), .CK(clk), .RN(n4447), .Q(
        \key_mem[3][82] ) );
  DFFRX1 \key_mem_reg[7][82]  ( .D(n2679), .CK(clk), .RN(n4447), .Q(
        \key_mem[7][82] ) );
  DFFRX1 \key_mem_reg[11][82]  ( .D(n3191), .CK(clk), .RN(n4448), .Q(
        \key_mem[11][82] ) );
  DFFRX1 \key_mem_reg[3][81]  ( .D(n2168), .CK(clk), .RN(n4449), .Q(
        \key_mem[3][81] ) );
  DFFRX1 \key_mem_reg[7][81]  ( .D(n2680), .CK(clk), .RN(n4449), .Q(
        \key_mem[7][81] ) );
  DFFRX1 \key_mem_reg[11][81]  ( .D(n3192), .CK(clk), .RN(n4450), .Q(
        \key_mem[11][81] ) );
  DFFRX1 \key_mem_reg[3][80]  ( .D(n2169), .CK(clk), .RN(n4450), .Q(
        \key_mem[3][80] ) );
  DFFRX1 \key_mem_reg[7][80]  ( .D(n2681), .CK(clk), .RN(n4451), .Q(
        \key_mem[7][80] ) );
  DFFRX1 \key_mem_reg[11][80]  ( .D(n3193), .CK(clk), .RN(n4451), .Q(
        \key_mem[11][80] ) );
  DFFRX1 \key_mem_reg[3][79]  ( .D(n2170), .CK(clk), .RN(n4452), .Q(
        \key_mem[3][79] ) );
  DFFRX1 \key_mem_reg[7][79]  ( .D(n2682), .CK(clk), .RN(n4453), .Q(
        \key_mem[7][79] ) );
  DFFRX1 \key_mem_reg[11][79]  ( .D(n3194), .CK(clk), .RN(n4453), .Q(
        \key_mem[11][79] ) );
  DFFRX1 \key_mem_reg[3][78]  ( .D(n2171), .CK(clk), .RN(n4454), .Q(
        \key_mem[3][78] ) );
  DFFRX1 \key_mem_reg[7][78]  ( .D(n2683), .CK(clk), .RN(n4454), .Q(
        \key_mem[7][78] ) );
  DFFRX1 \key_mem_reg[11][78]  ( .D(n3195), .CK(clk), .RN(n4455), .Q(
        \key_mem[11][78] ) );
  DFFRX1 \key_mem_reg[3][77]  ( .D(n2172), .CK(clk), .RN(n4388), .Q(
        \key_mem[3][77] ) );
  DFFRX1 \key_mem_reg[7][77]  ( .D(n2684), .CK(clk), .RN(n4373), .Q(
        \key_mem[7][77] ) );
  DFFRX1 \key_mem_reg[11][77]  ( .D(n3196), .CK(clk), .RN(n4374), .Q(
        \key_mem[11][77] ) );
  DFFRX1 \key_mem_reg[3][76]  ( .D(n2173), .CK(clk), .RN(n4374), .Q(
        \key_mem[3][76] ) );
  DFFRX1 \key_mem_reg[7][76]  ( .D(n2685), .CK(clk), .RN(n4375), .Q(
        \key_mem[7][76] ) );
  DFFRX1 \key_mem_reg[11][76]  ( .D(n3197), .CK(clk), .RN(n4375), .Q(
        \key_mem[11][76] ) );
  DFFRX1 \key_mem_reg[3][75]  ( .D(n2174), .CK(clk), .RN(n4376), .Q(
        \key_mem[3][75] ) );
  DFFRX1 \key_mem_reg[7][75]  ( .D(n2686), .CK(clk), .RN(n4377), .Q(
        \key_mem[7][75] ) );
  DFFRX1 \key_mem_reg[11][75]  ( .D(n3198), .CK(clk), .RN(n4377), .Q(
        \key_mem[11][75] ) );
  DFFRX1 \key_mem_reg[3][74]  ( .D(n2175), .CK(clk), .RN(n4378), .Q(
        \key_mem[3][74] ) );
  DFFRX1 \key_mem_reg[7][74]  ( .D(n2687), .CK(clk), .RN(n4378), .Q(
        \key_mem[7][74] ) );
  DFFRX1 \key_mem_reg[11][74]  ( .D(n3199), .CK(clk), .RN(n4379), .Q(
        \key_mem[11][74] ) );
  DFFRX1 \key_mem_reg[3][73]  ( .D(n2176), .CK(clk), .RN(n4380), .Q(
        \key_mem[3][73] ) );
  DFFRX1 \key_mem_reg[7][73]  ( .D(n2688), .CK(clk), .RN(n4380), .Q(
        \key_mem[7][73] ) );
  DFFRX1 \key_mem_reg[11][73]  ( .D(n3200), .CK(clk), .RN(n4381), .Q(
        \key_mem[11][73] ) );
  DFFRX1 \key_mem_reg[3][72]  ( .D(n2177), .CK(clk), .RN(n4381), .Q(
        \key_mem[3][72] ) );
  DFFRX1 \key_mem_reg[7][72]  ( .D(n2689), .CK(clk), .RN(n4382), .Q(
        \key_mem[7][72] ) );
  DFFRX1 \key_mem_reg[11][72]  ( .D(n3201), .CK(clk), .RN(n4382), .Q(
        \key_mem[11][72] ) );
  DFFRX1 \key_mem_reg[3][71]  ( .D(n2178), .CK(clk), .RN(n4383), .Q(
        \key_mem[3][71] ) );
  DFFRX1 \key_mem_reg[7][71]  ( .D(n2690), .CK(clk), .RN(n4384), .Q(
        \key_mem[7][71] ) );
  DFFRX1 \key_mem_reg[11][71]  ( .D(n3202), .CK(clk), .RN(n4384), .Q(
        \key_mem[11][71] ) );
  DFFRX1 \key_mem_reg[3][70]  ( .D(n2179), .CK(clk), .RN(n4385), .Q(
        \key_mem[3][70] ) );
  DFFRX1 \key_mem_reg[7][70]  ( .D(n2691), .CK(clk), .RN(n4385), .Q(
        \key_mem[7][70] ) );
  DFFRX1 \key_mem_reg[11][70]  ( .D(n3203), .CK(clk), .RN(n4386), .Q(
        \key_mem[11][70] ) );
  DFFRX1 \key_mem_reg[3][69]  ( .D(n2180), .CK(clk), .RN(n4387), .Q(
        \key_mem[3][69] ) );
  DFFRX1 \key_mem_reg[7][69]  ( .D(n2692), .CK(clk), .RN(n4387), .Q(
        \key_mem[7][69] ) );
  DFFRX1 \key_mem_reg[11][69]  ( .D(n3204), .CK(clk), .RN(n4388), .Q(
        \key_mem[11][69] ) );
  DFFRX1 \key_mem_reg[3][68]  ( .D(n2181), .CK(clk), .RN(n4558), .Q(
        \key_mem[3][68] ) );
  DFFRX1 \key_mem_reg[7][68]  ( .D(n2693), .CK(clk), .RN(n4381), .Q(
        \key_mem[7][68] ) );
  DFFRX1 \key_mem_reg[11][68]  ( .D(n3205), .CK(clk), .RN(n4401), .Q(
        \key_mem[11][68] ) );
  DFFRX1 \key_mem_reg[3][67]  ( .D(n2182), .CK(clk), .RN(n4389), .Q(
        \key_mem[3][67] ) );
  DFFRX1 \key_mem_reg[7][67]  ( .D(n2694), .CK(clk), .RN(n4379), .Q(
        \key_mem[7][67] ) );
  DFFRX1 \key_mem_reg[11][67]  ( .D(n3206), .CK(clk), .RN(n4378), .Q(
        \key_mem[11][67] ) );
  DFFRX1 \key_mem_reg[3][66]  ( .D(n2183), .CK(clk), .RN(n4399), .Q(
        \key_mem[3][66] ) );
  DFFRX1 \key_mem_reg[7][66]  ( .D(n2695), .CK(clk), .RN(n4398), .Q(
        \key_mem[7][66] ) );
  DFFRX1 \key_mem_reg[11][66]  ( .D(n3207), .CK(clk), .RN(n4461), .Q(
        \key_mem[11][66] ) );
  DFFRX1 \key_mem_reg[3][65]  ( .D(n2184), .CK(clk), .RN(n4455), .Q(
        \key_mem[3][65] ) );
  DFFRX1 \key_mem_reg[7][65]  ( .D(n2696), .CK(clk), .RN(n4456), .Q(
        \key_mem[7][65] ) );
  DFFRX1 \key_mem_reg[11][65]  ( .D(n3208), .CK(clk), .RN(n4447), .Q(
        \key_mem[11][65] ) );
  DFFRX1 \key_mem_reg[3][64]  ( .D(n2185), .CK(clk), .RN(n4448), .Q(
        \key_mem[3][64] ) );
  DFFRX1 \key_mem_reg[7][64]  ( .D(n2697), .CK(clk), .RN(n4422), .Q(
        \key_mem[7][64] ) );
  DFFRX1 \key_mem_reg[11][64]  ( .D(n3209), .CK(clk), .RN(n4419), .Q(
        \key_mem[11][64] ) );
  DFFRX1 \key_mem_reg[3][55]  ( .D(n2194), .CK(clk), .RN(n4513), .Q(
        \key_mem[3][55] ) );
  DFFRX1 \key_mem_reg[7][55]  ( .D(n2706), .CK(clk), .RN(n4547), .Q(
        \key_mem[7][55] ) );
  DFFRX1 \key_mem_reg[11][55]  ( .D(n3218), .CK(clk), .RN(n4546), .Q(
        \key_mem[11][55] ) );
  DFFRX1 \key_mem_reg[3][54]  ( .D(n2195), .CK(clk), .RN(n4542), .Q(
        \key_mem[3][54] ) );
  DFFRX1 \key_mem_reg[7][54]  ( .D(n2707), .CK(clk), .RN(n4541), .Q(
        \key_mem[7][54] ) );
  DFFRX1 \key_mem_reg[11][54]  ( .D(n3219), .CK(clk), .RN(n4370), .Q(
        \key_mem[11][54] ) );
  DFFRX1 \key_mem_reg[3][53]  ( .D(n2196), .CK(clk), .RN(n4371), .Q(
        \key_mem[3][53] ) );
  DFFRX1 \key_mem_reg[7][53]  ( .D(n2708), .CK(clk), .RN(n4371), .Q(
        \key_mem[7][53] ) );
  DFFRX1 \key_mem_reg[11][53]  ( .D(n3220), .CK(clk), .RN(n4372), .Q(
        \key_mem[11][53] ) );
  DFFRX1 \key_mem_reg[3][52]  ( .D(n2197), .CK(clk), .RN(n4372), .Q(
        \key_mem[3][52] ) );
  DFFRX1 \key_mem_reg[7][52]  ( .D(n2709), .CK(clk), .RN(n4403), .Q(
        \key_mem[7][52] ) );
  DFFRX1 \key_mem_reg[11][52]  ( .D(n3221), .CK(clk), .RN(n4404), .Q(
        \key_mem[11][52] ) );
  DFFRX1 \key_mem_reg[3][51]  ( .D(n2198), .CK(clk), .RN(n4404), .Q(
        \key_mem[3][51] ) );
  DFFRX1 \key_mem_reg[7][51]  ( .D(n2710), .CK(clk), .RN(n4405), .Q(
        \key_mem[7][51] ) );
  DFFRX1 \key_mem_reg[11][51]  ( .D(n3222), .CK(clk), .RN(n4405), .Q(
        \key_mem[11][51] ) );
  DFFRX1 \key_mem_reg[3][50]  ( .D(n2199), .CK(clk), .RN(n4406), .Q(
        \key_mem[3][50] ) );
  DFFRX1 \key_mem_reg[7][50]  ( .D(n2711), .CK(clk), .RN(n4407), .Q(
        \key_mem[7][50] ) );
  DFFRX1 \key_mem_reg[11][50]  ( .D(n3223), .CK(clk), .RN(n4407), .Q(
        \key_mem[11][50] ) );
  DFFRX1 \key_mem_reg[3][49]  ( .D(n2200), .CK(clk), .RN(n4408), .Q(
        \key_mem[3][49] ) );
  DFFRX1 \key_mem_reg[7][49]  ( .D(n2712), .CK(clk), .RN(n4408), .Q(
        \key_mem[7][49] ) );
  DFFRX1 \key_mem_reg[11][49]  ( .D(n3224), .CK(clk), .RN(n4409), .Q(
        \key_mem[11][49] ) );
  DFFRX1 \key_mem_reg[3][47]  ( .D(n2202), .CK(clk), .RN(n4411), .Q(
        \key_mem[3][47] ) );
  DFFRX1 \key_mem_reg[7][47]  ( .D(n2714), .CK(clk), .RN(n4412), .Q(
        \key_mem[7][47] ) );
  DFFRX1 \key_mem_reg[11][47]  ( .D(n3226), .CK(clk), .RN(n4412), .Q(
        \key_mem[11][47] ) );
  DFFRX1 \key_mem_reg[3][46]  ( .D(n2203), .CK(clk), .RN(n4413), .Q(
        \key_mem[3][46] ) );
  DFFRX1 \key_mem_reg[7][46]  ( .D(n2715), .CK(clk), .RN(n4411), .Q(
        \key_mem[7][46] ) );
  DFFRX1 \key_mem_reg[11][46]  ( .D(n3227), .CK(clk), .RN(n4410), .Q(
        \key_mem[11][46] ) );
  DFFRX1 \key_mem_reg[3][45]  ( .D(n2204), .CK(clk), .RN(n4414), .Q(
        \key_mem[3][45] ) );
  DFFRX1 \key_mem_reg[7][45]  ( .D(n2716), .CK(clk), .RN(n4414), .Q(
        \key_mem[7][45] ) );
  DFFRX1 \key_mem_reg[11][45]  ( .D(n3228), .CK(clk), .RN(n4415), .Q(
        \key_mem[11][45] ) );
  DFFRX1 \key_mem_reg[3][44]  ( .D(n2205), .CK(clk), .RN(n4416), .Q(
        \key_mem[3][44] ) );
  DFFRX1 \key_mem_reg[7][44]  ( .D(n2717), .CK(clk), .RN(n4416), .Q(
        \key_mem[7][44] ) );
  DFFRX1 \key_mem_reg[11][44]  ( .D(n3229), .CK(clk), .RN(n4417), .Q(
        \key_mem[11][44] ) );
  DFFRX1 \key_mem_reg[3][43]  ( .D(n2206), .CK(clk), .RN(n4388), .Q(
        \key_mem[3][43] ) );
  DFFRX1 \key_mem_reg[7][43]  ( .D(n2718), .CK(clk), .RN(n4389), .Q(
        \key_mem[7][43] ) );
  DFFRX1 \key_mem_reg[11][43]  ( .D(n3230), .CK(clk), .RN(n4389), .Q(
        \key_mem[11][43] ) );
  DFFRX1 \key_mem_reg[3][42]  ( .D(n2207), .CK(clk), .RN(n4390), .Q(
        \key_mem[3][42] ) );
  DFFRX1 \key_mem_reg[7][42]  ( .D(n2719), .CK(clk), .RN(n4390), .Q(
        \key_mem[7][42] ) );
  DFFRX1 \key_mem_reg[11][42]  ( .D(n3231), .CK(clk), .RN(n4391), .Q(
        \key_mem[11][42] ) );
  DFFRX1 \key_mem_reg[3][41]  ( .D(n2208), .CK(clk), .RN(n4392), .Q(
        \key_mem[3][41] ) );
  DFFRX1 \key_mem_reg[7][41]  ( .D(n2720), .CK(clk), .RN(n4392), .Q(
        \key_mem[7][41] ) );
  DFFRX1 \key_mem_reg[11][41]  ( .D(n3232), .CK(clk), .RN(n4393), .Q(
        \key_mem[11][41] ) );
  DFFRX1 \key_mem_reg[3][40]  ( .D(n2209), .CK(clk), .RN(n4393), .Q(
        \key_mem[3][40] ) );
  DFFRX1 \key_mem_reg[7][40]  ( .D(n2721), .CK(clk), .RN(n4394), .Q(
        \key_mem[7][40] ) );
  DFFRX1 \key_mem_reg[11][40]  ( .D(n3233), .CK(clk), .RN(n4394), .Q(
        \key_mem[11][40] ) );
  DFFRX1 \key_mem_reg[3][39]  ( .D(n2210), .CK(clk), .RN(n4395), .Q(
        \key_mem[3][39] ) );
  DFFRX1 \key_mem_reg[7][39]  ( .D(n2722), .CK(clk), .RN(n4396), .Q(
        \key_mem[7][39] ) );
  DFFRX1 \key_mem_reg[11][39]  ( .D(n3234), .CK(clk), .RN(n4396), .Q(
        \key_mem[11][39] ) );
  DFFRX1 \key_mem_reg[3][38]  ( .D(n2211), .CK(clk), .RN(n4397), .Q(
        \key_mem[3][38] ) );
  DFFRX1 \key_mem_reg[7][38]  ( .D(n2723), .CK(clk), .RN(n4398), .Q(
        \key_mem[7][38] ) );
  DFFRX1 \key_mem_reg[11][38]  ( .D(n3235), .CK(clk), .RN(n4398), .Q(
        \key_mem[11][38] ) );
  DFFRX1 \key_mem_reg[3][37]  ( .D(n2212), .CK(clk), .RN(n4399), .Q(
        \key_mem[3][37] ) );
  DFFRX1 \key_mem_reg[7][37]  ( .D(n2724), .CK(clk), .RN(n4399), .Q(
        \key_mem[7][37] ) );
  DFFRX1 \key_mem_reg[11][37]  ( .D(n3236), .CK(clk), .RN(n4400), .Q(
        \key_mem[11][37] ) );
  DFFRX1 \key_mem_reg[3][36]  ( .D(n2213), .CK(clk), .RN(n4401), .Q(
        \key_mem[3][36] ) );
  DFFRX1 \key_mem_reg[7][36]  ( .D(n2725), .CK(clk), .RN(n4401), .Q(
        \key_mem[7][36] ) );
  DFFRX1 \key_mem_reg[11][36]  ( .D(n3237), .CK(clk), .RN(n4402), .Q(
        \key_mem[11][36] ) );
  DFFRX1 \key_mem_reg[3][35]  ( .D(n2214), .CK(clk), .RN(n4402), .Q(
        \key_mem[3][35] ) );
  DFFRX1 \key_mem_reg[7][35]  ( .D(n2726), .CK(clk), .RN(n4403), .Q(
        \key_mem[7][35] ) );
  DFFRX1 \key_mem_reg[11][35]  ( .D(n3238), .CK(clk), .RN(n4549), .Q(
        \key_mem[11][35] ) );
  DFFRX1 \key_mem_reg[3][34]  ( .D(n2215), .CK(clk), .RN(n4542), .Q(
        \key_mem[3][34] ) );
  DFFRX1 \key_mem_reg[7][34]  ( .D(n2727), .CK(clk), .RN(n4542), .Q(
        \key_mem[7][34] ) );
  DFFRX1 \key_mem_reg[11][34]  ( .D(n3239), .CK(clk), .RN(n4543), .Q(
        \key_mem[11][34] ) );
  DFFRX1 \key_mem_reg[3][33]  ( .D(n2216), .CK(clk), .RN(n4544), .Q(
        \key_mem[3][33] ) );
  DFFRX1 \key_mem_reg[7][33]  ( .D(n2728), .CK(clk), .RN(n4544), .Q(
        \key_mem[7][33] ) );
  DFFRX1 \key_mem_reg[11][33]  ( .D(n3240), .CK(clk), .RN(n4545), .Q(
        \key_mem[11][33] ) );
  DFFRX1 \key_mem_reg[3][32]  ( .D(n2217), .CK(clk), .RN(n4545), .Q(
        \key_mem[3][32] ) );
  DFFRX1 \key_mem_reg[7][32]  ( .D(n2729), .CK(clk), .RN(n4546), .Q(
        \key_mem[7][32] ) );
  DFFRX1 \key_mem_reg[11][32]  ( .D(n3241), .CK(clk), .RN(n4546), .Q(
        \key_mem[11][32] ) );
  DFFRX1 \key_mem_reg[3][23]  ( .D(n2226), .CK(clk), .RN(n4547), .Q(
        \key_mem[3][23] ) );
  DFFRX1 \key_mem_reg[7][23]  ( .D(n2738), .CK(clk), .RN(n4548), .Q(
        \key_mem[7][23] ) );
  DFFRX1 \key_mem_reg[11][23]  ( .D(n3250), .CK(clk), .RN(n4548), .Q(
        \key_mem[11][23] ) );
  DFFRX1 \key_mem_reg[3][22]  ( .D(n2227), .CK(clk), .RN(n4549), .Q(
        \key_mem[3][22] ) );
  DFFRX1 \key_mem_reg[7][22]  ( .D(n2739), .CK(clk), .RN(n4550), .Q(
        \key_mem[7][22] ) );
  DFFRX1 \key_mem_reg[11][22]  ( .D(n3251), .CK(clk), .RN(n4550), .Q(
        \key_mem[11][22] ) );
  DFFRX1 \key_mem_reg[3][21]  ( .D(n2228), .CK(clk), .RN(n4551), .Q(
        \key_mem[3][21] ) );
  DFFRX1 \key_mem_reg[7][21]  ( .D(n2740), .CK(clk), .RN(n4551), .Q(
        \key_mem[7][21] ) );
  DFFRX1 \key_mem_reg[11][21]  ( .D(n3252), .CK(clk), .RN(n4552), .Q(
        \key_mem[11][21] ) );
  DFFRX1 \key_mem_reg[3][20]  ( .D(n2229), .CK(clk), .RN(n4553), .Q(
        \key_mem[3][20] ) );
  DFFRX1 \key_mem_reg[7][20]  ( .D(n2741), .CK(clk), .RN(n4553), .Q(
        \key_mem[7][20] ) );
  DFFRX1 \key_mem_reg[11][20]  ( .D(n3253), .CK(clk), .RN(n4424), .Q(
        \key_mem[11][20] ) );
  DFFRX1 \key_mem_reg[3][18]  ( .D(n2231), .CK(clk), .RN(n4554), .Q(
        \key_mem[3][18] ) );
  DFFRX1 \key_mem_reg[7][18]  ( .D(n2743), .CK(clk), .RN(n4526), .Q(
        \key_mem[7][18] ) );
  DFFRX1 \key_mem_reg[11][18]  ( .D(n3255), .CK(clk), .RN(n4527), .Q(
        \key_mem[11][18] ) );
  DFFRX1 \key_mem_reg[3][16]  ( .D(n2233), .CK(clk), .RN(n4529), .Q(
        \key_mem[3][16] ) );
  DFFRX1 \key_mem_reg[7][16]  ( .D(n2745), .CK(clk), .RN(n4530), .Q(
        \key_mem[7][16] ) );
  DFFRX1 \key_mem_reg[11][16]  ( .D(n3257), .CK(clk), .RN(n4530), .Q(
        \key_mem[11][16] ) );
  DFFRX1 \key_mem_reg[3][15]  ( .D(n2234), .CK(clk), .RN(n4531), .Q(
        \key_mem[3][15] ) );
  DFFRX1 \key_mem_reg[7][15]  ( .D(n2746), .CK(clk), .RN(n4532), .Q(
        \key_mem[7][15] ) );
  DFFRX1 \key_mem_reg[11][15]  ( .D(n3258), .CK(clk), .RN(n4532), .Q(
        \key_mem[11][15] ) );
  DFFRX1 \key_mem_reg[3][14]  ( .D(n2235), .CK(clk), .RN(n4533), .Q(
        \key_mem[3][14] ) );
  DFFRX1 \key_mem_reg[7][14]  ( .D(n2747), .CK(clk), .RN(n4533), .Q(
        \key_mem[7][14] ) );
  DFFRX1 \key_mem_reg[11][14]  ( .D(n3259), .CK(clk), .RN(n4534), .Q(
        \key_mem[11][14] ) );
  DFFRX1 \key_mem_reg[3][13]  ( .D(n2236), .CK(clk), .RN(n4535), .Q(
        \key_mem[3][13] ) );
  DFFRX1 \key_mem_reg[7][13]  ( .D(n2748), .CK(clk), .RN(n4535), .Q(
        \key_mem[7][13] ) );
  DFFRX1 \key_mem_reg[11][13]  ( .D(n3260), .CK(clk), .RN(n4536), .Q(
        \key_mem[11][13] ) );
  DFFRX1 \key_mem_reg[3][12]  ( .D(n2237), .CK(clk), .RN(n4536), .Q(
        \key_mem[3][12] ) );
  DFFRX1 \key_mem_reg[7][12]  ( .D(n2749), .CK(clk), .RN(n4537), .Q(
        \key_mem[7][12] ) );
  DFFRX1 \key_mem_reg[11][12]  ( .D(n3261), .CK(clk), .RN(n4537), .Q(
        \key_mem[11][12] ) );
  DFFRX1 \key_mem_reg[3][11]  ( .D(n2238), .CK(clk), .RN(n4538), .Q(
        \key_mem[3][11] ) );
  DFFRX1 \key_mem_reg[7][11]  ( .D(n2750), .CK(clk), .RN(n4539), .Q(
        \key_mem[7][11] ) );
  DFFRX1 \key_mem_reg[11][11]  ( .D(n3262), .CK(clk), .RN(n4539), .Q(
        \key_mem[11][11] ) );
  DFFRX1 \key_mem_reg[3][10]  ( .D(n2239), .CK(clk), .RN(n4540), .Q(
        \key_mem[3][10] ) );
  DFFRX1 \key_mem_reg[7][10]  ( .D(n2751), .CK(clk), .RN(n4540), .Q(
        \key_mem[7][10] ) );
  DFFRX1 \key_mem_reg[11][10]  ( .D(n3263), .CK(clk), .RN(n4541), .Q(
        \key_mem[11][10] ) );
  DFFRX1 \key_mem_reg[3][9]  ( .D(n2240), .CK(clk), .RN(n4535), .Q(
        \key_mem[3][9] ) );
  DFFRX1 \key_mem_reg[7][9]  ( .D(n2752), .CK(clk), .RN(n4534), .Q(
        \key_mem[7][9] ) );
  DFFRX1 \key_mem_reg[11][9]  ( .D(n3264), .CK(clk), .RN(n4530), .Q(
        \key_mem[11][9] ) );
  DFFRX1 \key_mem_reg[3][8]  ( .D(n2241), .CK(clk), .RN(n4496), .Q(
        \key_mem[3][8] ) );
  DFFRX1 \key_mem_reg[7][8]  ( .D(n2753), .CK(clk), .RN(n4494), .Q(
        \key_mem[7][8] ) );
  DFFRX1 \key_mem_reg[11][8]  ( .D(n3265), .CK(clk), .RN(n4559), .Q(
        \key_mem[11][8] ) );
  DFFRX1 \key_mem_reg[3][7]  ( .D(n2242), .CK(clk), .RN(n4559), .Q(
        \key_mem[3][7] ) );
  DFFRX1 \key_mem_reg[7][7]  ( .D(n2754), .CK(clk), .RN(n4560), .Q(
        \key_mem[7][7] ) );
  DFFRX1 \key_mem_reg[11][7]  ( .D(n3266), .CK(clk), .RN(n4560), .Q(
        \key_mem[11][7] ) );
  DFFRX1 \key_mem_reg[3][6]  ( .D(n2243), .CK(clk), .RN(n4561), .Q(
        \key_mem[3][6] ) );
  DFFRX1 \key_mem_reg[7][6]  ( .D(n2755), .CK(clk), .RN(n4562), .Q(
        \key_mem[7][6] ) );
  DFFRX1 \key_mem_reg[11][6]  ( .D(n3267), .CK(clk), .RN(n4562), .Q(
        \key_mem[11][6] ) );
  DFFRX1 \key_mem_reg[3][5]  ( .D(n2244), .CK(clk), .RN(n4374), .Q(
        \key_mem[3][5] ) );
  DFFRX1 \key_mem_reg[7][5]  ( .D(n2756), .CK(clk), .RN(n4442), .Q(
        \key_mem[7][5] ) );
  DFFRX1 \key_mem_reg[11][5]  ( .D(n3268), .CK(clk), .RN(n4432), .Q(
        \key_mem[11][5] ) );
  DFFRX1 \key_mem_reg[3][4]  ( .D(n2245), .CK(clk), .RN(n4411), .Q(
        \key_mem[3][4] ) );
  DFFRX1 \key_mem_reg[7][4]  ( .D(n2757), .CK(clk), .RN(n4410), .Q(
        \key_mem[7][4] ) );
  DFFRX1 \key_mem_reg[11][4]  ( .D(n3269), .CK(clk), .RN(n4464), .Q(
        \key_mem[11][4] ) );
  DFFRX1 \key_mem_reg[3][3]  ( .D(n2246), .CK(clk), .RN(n4389), .Q(
        \key_mem[3][3] ) );
  DFFRX1 \key_mem_reg[7][3]  ( .D(n2758), .CK(clk), .RN(n4379), .Q(
        \key_mem[7][3] ) );
  DFFRX1 \key_mem_reg[11][3]  ( .D(n3270), .CK(clk), .RN(n4384), .Q(
        \key_mem[11][3] ) );
  DFFRX1 \key_mem_reg[3][2]  ( .D(n2247), .CK(clk), .RN(n4417), .Q(
        \key_mem[3][2] ) );
  DFFRX1 \key_mem_reg[7][2]  ( .D(n2759), .CK(clk), .RN(n4563), .Q(
        \key_mem[7][2] ) );
  DFFRX1 \key_mem_reg[11][2]  ( .D(n3271), .CK(clk), .RN(n4563), .Q(
        \key_mem[11][2] ) );
  DFFRX1 \key_mem_reg[3][1]  ( .D(n2248), .CK(clk), .RN(n4564), .Q(
        \key_mem[3][1] ) );
  DFFRX1 \key_mem_reg[7][1]  ( .D(n2760), .CK(clk), .RN(n4564), .Q(
        \key_mem[7][1] ) );
  DFFRX1 \key_mem_reg[11][1]  ( .D(n3272), .CK(clk), .RN(n4555), .Q(
        \key_mem[11][1] ) );
  DFFRX1 \key_mem_reg[3][0]  ( .D(n2249), .CK(clk), .RN(n4555), .Q(
        \key_mem[3][0] ) );
  DFFRX1 \key_mem_reg[7][0]  ( .D(n2761), .CK(clk), .RN(n4556), .Q(
        \key_mem[7][0] ) );
  DFFRX1 \key_mem_reg[11][0]  ( .D(n3273), .CK(clk), .RN(n4556), .Q(
        \key_mem[11][0] ) );
  DFFRX1 \key_mem_reg[3][127]  ( .D(n2122), .CK(clk), .RN(n4490), .Q(
        \key_mem[3][127] ) );
  DFFRX1 \key_mem_reg[7][127]  ( .D(n2634), .CK(clk), .RN(n4533), .Q(
        \key_mem[7][127] ) );
  DFFRX1 \key_mem_reg[11][127]  ( .D(n3146), .CK(clk), .RN(n4532), .Q(
        \key_mem[11][127] ) );
  DFFRX1 \key_mem_reg[3][95]  ( .D(n2154), .CK(clk), .RN(n4524), .Q(
        \key_mem[3][95] ) );
  DFFRX1 \key_mem_reg[7][95]  ( .D(n2666), .CK(clk), .RN(n4514), .Q(
        \key_mem[7][95] ) );
  DFFRX1 \key_mem_reg[11][95]  ( .D(n3178), .CK(clk), .RN(n4513), .Q(
        \key_mem[11][95] ) );
  DFFRX1 \key_mem_reg[3][63]  ( .D(n2186), .CK(clk), .RN(n4562), .Q(
        \key_mem[3][63] ) );
  DFFRX1 \key_mem_reg[7][63]  ( .D(n2698), .CK(clk), .RN(n4561), .Q(
        \key_mem[7][63] ) );
  DFFRX1 \key_mem_reg[11][63]  ( .D(n3210), .CK(clk), .RN(n4558), .Q(
        \key_mem[11][63] ) );
  DFFRX1 \key_mem_reg[3][31]  ( .D(n2218), .CK(clk), .RN(n4557), .Q(
        \key_mem[3][31] ) );
  DFFRX1 \key_mem_reg[7][31]  ( .D(n2730), .CK(clk), .RN(n4557), .Q(
        \key_mem[7][31] ) );
  DFFRX1 \key_mem_reg[11][31]  ( .D(n3242), .CK(clk), .RN(n4459), .Q(
        \key_mem[11][31] ) );
  DFFRX1 \key_mem_reg[3][120]  ( .D(n2129), .CK(clk), .RN(n4491), .Q(
        \key_mem[3][120] ) );
  DFFRX1 \key_mem_reg[7][120]  ( .D(n2641), .CK(clk), .RN(n4490), .Q(
        \key_mem[7][120] ) );
  DFFRX1 \key_mem_reg[11][120]  ( .D(n3153), .CK(clk), .RN(n4547), .Q(
        \key_mem[11][120] ) );
  DFFRX1 \key_mem_reg[3][88]  ( .D(n2161), .CK(clk), .RN(n4546), .Q(
        \key_mem[3][88] ) );
  DFFRX1 \key_mem_reg[7][88]  ( .D(n2673), .CK(clk), .RN(n4558), .Q(
        \key_mem[7][88] ) );
  DFFRX1 \key_mem_reg[11][88]  ( .D(n3185), .CK(clk), .RN(n4558), .Q(
        \key_mem[11][88] ) );
  DFFRX1 \key_mem_reg[3][56]  ( .D(n2193), .CK(clk), .RN(n4475), .Q(
        \key_mem[3][56] ) );
  DFFRX1 \key_mem_reg[7][56]  ( .D(n2705), .CK(clk), .RN(n4511), .Q(
        \key_mem[7][56] ) );
  DFFRX1 \key_mem_reg[11][56]  ( .D(n3217), .CK(clk), .RN(n4510), .Q(
        \key_mem[11][56] ) );
  DFFRX1 \key_mem_reg[3][24]  ( .D(n2225), .CK(clk), .RN(n4451), .Q(
        \key_mem[3][24] ) );
  DFFRX1 \key_mem_reg[7][24]  ( .D(n2737), .CK(clk), .RN(n4452), .Q(
        \key_mem[7][24] ) );
  DFFRX1 \key_mem_reg[11][24]  ( .D(n3249), .CK(clk), .RN(n4553), .Q(
        \key_mem[11][24] ) );
  DFFRX1 \key_mem_reg[3][122]  ( .D(n2127), .CK(clk), .RN(n4485), .Q(
        \key_mem[3][122] ) );
  DFFRX1 \key_mem_reg[7][122]  ( .D(n2639), .CK(clk), .RN(n4485), .Q(
        \key_mem[7][122] ) );
  DFFRX1 \key_mem_reg[11][122]  ( .D(n3151), .CK(clk), .RN(n4486), .Q(
        \key_mem[11][122] ) );
  DFFRX1 \key_mem_reg[3][90]  ( .D(n2159), .CK(clk), .RN(n4487), .Q(
        \key_mem[3][90] ) );
  DFFRX1 \key_mem_reg[7][90]  ( .D(n2671), .CK(clk), .RN(n4487), .Q(
        \key_mem[7][90] ) );
  DFFRX1 \key_mem_reg[11][90]  ( .D(n3183), .CK(clk), .RN(n4488), .Q(
        \key_mem[11][90] ) );
  DFFRX1 \key_mem_reg[3][58]  ( .D(n2191), .CK(clk), .RN(n4488), .Q(
        \key_mem[3][58] ) );
  DFFRX1 \key_mem_reg[7][58]  ( .D(n2703), .CK(clk), .RN(n4489), .Q(
        \key_mem[7][58] ) );
  DFFRX1 \key_mem_reg[11][58]  ( .D(n3215), .CK(clk), .RN(n4489), .Q(
        \key_mem[11][58] ) );
  DFFRX1 \key_mem_reg[3][26]  ( .D(n2223), .CK(clk), .RN(n4490), .Q(
        \key_mem[3][26] ) );
  DFFRX1 \key_mem_reg[7][26]  ( .D(n2735), .CK(clk), .RN(n4491), .Q(
        \key_mem[7][26] ) );
  DFFRX1 \key_mem_reg[11][26]  ( .D(n3247), .CK(clk), .RN(n4491), .Q(
        \key_mem[11][26] ) );
  DFFRX1 \key_mem_reg[3][123]  ( .D(n2126), .CK(clk), .RN(n4557), .Q(
        \key_mem[3][123] ) );
  DFFRX1 \key_mem_reg[7][123]  ( .D(n2638), .CK(clk), .RN(n4431), .Q(
        \key_mem[7][123] ) );
  DFFRX1 \key_mem_reg[11][123]  ( .D(n3150), .CK(clk), .RN(n4432), .Q(
        \key_mem[11][123] ) );
  DFFRX1 \key_mem_reg[3][91]  ( .D(n2158), .CK(clk), .RN(n4492), .Q(
        \key_mem[3][91] ) );
  DFFRX1 \key_mem_reg[7][91]  ( .D(n2670), .CK(clk), .RN(n4492), .Q(
        \key_mem[7][91] ) );
  DFFRX1 \key_mem_reg[11][91]  ( .D(n3182), .CK(clk), .RN(n4493), .Q(
        \key_mem[11][91] ) );
  DFFRX1 \key_mem_reg[3][59]  ( .D(n2190), .CK(clk), .RN(n4494), .Q(
        \key_mem[3][59] ) );
  DFFRX1 \key_mem_reg[7][59]  ( .D(n2702), .CK(clk), .RN(n4494), .Q(
        \key_mem[7][59] ) );
  DFFRX1 \key_mem_reg[11][59]  ( .D(n3214), .CK(clk), .RN(n4495), .Q(
        \key_mem[11][59] ) );
  DFFRX1 \key_mem_reg[3][27]  ( .D(n2222), .CK(clk), .RN(n4495), .Q(
        \key_mem[3][27] ) );
  DFFRX1 \key_mem_reg[7][27]  ( .D(n2734), .CK(clk), .RN(n4477), .Q(
        \key_mem[7][27] ) );
  DFFRX1 \key_mem_reg[11][27]  ( .D(n3246), .CK(clk), .RN(n4470), .Q(
        \key_mem[11][27] ) );
  DFFRX1 \key_mem_reg[3][126]  ( .D(n2123), .CK(clk), .RN(n4471), .Q(
        \key_mem[3][126] ) );
  DFFRX1 \key_mem_reg[7][126]  ( .D(n2635), .CK(clk), .RN(n4472), .Q(
        \key_mem[7][126] ) );
  DFFRX1 \key_mem_reg[11][126]  ( .D(n3147), .CK(clk), .RN(n4472), .Q(
        \key_mem[11][126] ) );
  DFFRX1 \key_mem_reg[3][94]  ( .D(n2155), .CK(clk), .RN(n4473), .Q(
        \key_mem[3][94] ) );
  DFFRX1 \key_mem_reg[7][94]  ( .D(n2667), .CK(clk), .RN(n4473), .Q(
        \key_mem[7][94] ) );
  DFFRX1 \key_mem_reg[11][94]  ( .D(n3179), .CK(clk), .RN(n4474), .Q(
        \key_mem[11][94] ) );
  DFFRX1 \key_mem_reg[3][62]  ( .D(n2187), .CK(clk), .RN(n4475), .Q(
        \key_mem[3][62] ) );
  DFFRX1 \key_mem_reg[7][62]  ( .D(n2699), .CK(clk), .RN(n4475), .Q(
        \key_mem[7][62] ) );
  DFFRX1 \key_mem_reg[11][62]  ( .D(n3211), .CK(clk), .RN(n4476), .Q(
        \key_mem[11][62] ) );
  DFFRX1 \key_mem_reg[3][30]  ( .D(n2219), .CK(clk), .RN(n4476), .Q(
        \key_mem[3][30] ) );
  DFFRX1 \key_mem_reg[7][30]  ( .D(n2731), .CK(clk), .RN(n4477), .Q(
        \key_mem[7][30] ) );
  DFFRX1 \key_mem_reg[11][30]  ( .D(n3243), .CK(clk), .RN(n4478), .Q(
        \key_mem[11][30] ) );
  DFFRX1 \key_mem_reg[3][125]  ( .D(n2124), .CK(clk), .RN(n4478), .Q(
        \key_mem[3][125] ) );
  DFFRX1 \key_mem_reg[7][125]  ( .D(n2636), .CK(clk), .RN(n4479), .Q(
        \key_mem[7][125] ) );
  DFFRX1 \key_mem_reg[11][125]  ( .D(n3148), .CK(clk), .RN(n4479), .Q(
        \key_mem[11][125] ) );
  DFFRX1 \key_mem_reg[3][93]  ( .D(n2156), .CK(clk), .RN(n4480), .Q(
        \key_mem[3][93] ) );
  DFFRX1 \key_mem_reg[7][93]  ( .D(n2668), .CK(clk), .RN(n4481), .Q(
        \key_mem[7][93] ) );
  DFFRX1 \key_mem_reg[11][93]  ( .D(n3180), .CK(clk), .RN(n4481), .Q(
        \key_mem[11][93] ) );
  DFFRX1 \key_mem_reg[3][61]  ( .D(n2188), .CK(clk), .RN(n4482), .Q(
        \key_mem[3][61] ) );
  DFFRX1 \key_mem_reg[7][61]  ( .D(n2700), .CK(clk), .RN(n4482), .Q(
        \key_mem[7][61] ) );
  DFFRX1 \key_mem_reg[11][61]  ( .D(n3212), .CK(clk), .RN(n4483), .Q(
        \key_mem[11][61] ) );
  DFFRX1 \key_mem_reg[3][29]  ( .D(n2220), .CK(clk), .RN(n4484), .Q(
        \key_mem[3][29] ) );
  DFFRX1 \key_mem_reg[7][29]  ( .D(n2732), .CK(clk), .RN(n4484), .Q(
        \key_mem[7][29] ) );
  DFFRX1 \key_mem_reg[11][29]  ( .D(n3244), .CK(clk), .RN(n4449), .Q(
        \key_mem[11][29] ) );
  DFFRX1 \key_mem_reg[3][124]  ( .D(n2125), .CK(clk), .RN(n4511), .Q(
        \key_mem[3][124] ) );
  DFFRX1 \key_mem_reg[7][124]  ( .D(n2637), .CK(clk), .RN(n4512), .Q(
        \key_mem[7][124] ) );
  DFFRX1 \key_mem_reg[11][124]  ( .D(n3149), .CK(clk), .RN(n4512), .Q(
        \key_mem[11][124] ) );
  DFFRX1 \key_mem_reg[3][92]  ( .D(n2157), .CK(clk), .RN(n4513), .Q(
        \key_mem[3][92] ) );
  DFFRX1 \key_mem_reg[7][92]  ( .D(n2669), .CK(clk), .RN(n4514), .Q(
        \key_mem[7][92] ) );
  DFFRX1 \key_mem_reg[11][92]  ( .D(n3181), .CK(clk), .RN(n4514), .Q(
        \key_mem[11][92] ) );
  DFFRX1 \key_mem_reg[3][60]  ( .D(n2189), .CK(clk), .RN(n4515), .Q(
        \key_mem[3][60] ) );
  DFFRX1 \key_mem_reg[7][60]  ( .D(n2701), .CK(clk), .RN(n4515), .Q(
        \key_mem[7][60] ) );
  DFFRX1 \key_mem_reg[11][60]  ( .D(n3213), .CK(clk), .RN(n4516), .Q(
        \key_mem[11][60] ) );
  DFFRX1 \key_mem_reg[3][28]  ( .D(n2221), .CK(clk), .RN(n4517), .Q(
        \key_mem[3][28] ) );
  DFFRX1 \key_mem_reg[7][28]  ( .D(n2733), .CK(clk), .RN(n4517), .Q(
        \key_mem[7][28] ) );
  DFFRX1 \key_mem_reg[11][28]  ( .D(n3245), .CK(clk), .RN(n4518), .Q(
        \key_mem[11][28] ) );
  DFFRX1 \key_mem_reg[3][121]  ( .D(n2128), .CK(clk), .RN(n4519), .Q(
        \key_mem[3][121] ) );
  DFFRX1 \key_mem_reg[7][121]  ( .D(n2640), .CK(clk), .RN(n4519), .Q(
        \key_mem[7][121] ) );
  DFFRX1 \key_mem_reg[11][121]  ( .D(n3152), .CK(clk), .RN(n4520), .Q(
        \key_mem[11][121] ) );
  DFFRX1 \key_mem_reg[3][89]  ( .D(n2160), .CK(clk), .RN(n4520), .Q(
        \key_mem[3][89] ) );
  DFFRX1 \key_mem_reg[7][89]  ( .D(n2672), .CK(clk), .RN(n4521), .Q(
        \key_mem[7][89] ) );
  DFFRX1 \key_mem_reg[11][89]  ( .D(n3184), .CK(clk), .RN(n4521), .Q(
        \key_mem[11][89] ) );
  DFFRX1 \key_mem_reg[3][57]  ( .D(n2192), .CK(clk), .RN(n4522), .Q(
        \key_mem[3][57] ) );
  DFFRX1 \key_mem_reg[7][57]  ( .D(n2704), .CK(clk), .RN(n4523), .Q(
        \key_mem[7][57] ) );
  DFFRX1 \key_mem_reg[11][57]  ( .D(n3216), .CK(clk), .RN(n4523), .Q(
        \key_mem[11][57] ) );
  DFFRX1 \key_mem_reg[3][25]  ( .D(n2224), .CK(clk), .RN(n4524), .Q(
        \key_mem[3][25] ) );
  DFFRX1 \key_mem_reg[7][25]  ( .D(n2736), .CK(clk), .RN(n4524), .Q(
        \key_mem[7][25] ) );
  DFFRX1 \key_mem_reg[11][25]  ( .D(n3248), .CK(clk), .RN(n4525), .Q(
        \key_mem[11][25] ) );
  DFFRX1 \key_mem_reg[0][119]  ( .D(n1746), .CK(clk), .RN(n4430), .Q(
        \key_mem[0][119] ) );
  DFFRX1 \key_mem_reg[4][119]  ( .D(n2258), .CK(clk), .RN(n4430), .Q(
        \key_mem[4][119] ) );
  DFFRX1 \key_mem_reg[8][119]  ( .D(n2770), .CK(clk), .RN(n4431), .Q(
        \key_mem[8][119] ) );
  DFFRX1 \key_mem_reg[0][118]  ( .D(n1747), .CK(clk), .RN(n4431), .Q(
        \key_mem[0][118] ) );
  DFFRX1 \key_mem_reg[4][118]  ( .D(n2259), .CK(clk), .RN(n4432), .Q(
        \key_mem[4][118] ) );
  DFFRX1 \key_mem_reg[8][118]  ( .D(n2771), .CK(clk), .RN(n4432), .Q(
        \key_mem[8][118] ) );
  DFFRX1 \key_mem_reg[0][117]  ( .D(n1748), .CK(clk), .RN(n4371), .Q(
        \key_mem[0][117] ) );
  DFFRX1 \key_mem_reg[4][117]  ( .D(n2260), .CK(clk), .RN(n4433), .Q(
        \key_mem[4][117] ) );
  DFFRX1 \key_mem_reg[8][117]  ( .D(n2772), .CK(clk), .RN(n4433), .Q(
        \key_mem[8][117] ) );
  DFFRX1 \key_mem_reg[0][116]  ( .D(n1749), .CK(clk), .RN(n4497), .Q(
        \key_mem[0][116] ) );
  DFFRX1 \key_mem_reg[4][116]  ( .D(n2261), .CK(clk), .RN(n4496), .Q(
        \key_mem[4][116] ) );
  DFFRX1 \key_mem_reg[8][116]  ( .D(n2773), .CK(clk), .RN(n4402), .Q(
        \key_mem[8][116] ) );
  DFFRX1 \key_mem_reg[0][115]  ( .D(n1750), .CK(clk), .RN(n4395), .Q(
        \key_mem[0][115] ) );
  DFFRX1 \key_mem_reg[4][115]  ( .D(n2262), .CK(clk), .RN(n4394), .Q(
        \key_mem[4][115] ) );
  DFFRX1 \key_mem_reg[8][115]  ( .D(n2774), .CK(clk), .RN(n4434), .Q(
        \key_mem[8][115] ) );
  DFFRX1 \key_mem_reg[0][114]  ( .D(n1751), .CK(clk), .RN(n4435), .Q(
        \key_mem[0][114] ) );
  DFFRX1 \key_mem_reg[4][114]  ( .D(n2263), .CK(clk), .RN(n4435), .Q(
        \key_mem[4][114] ) );
  DFFRX1 \key_mem_reg[8][114]  ( .D(n2775), .CK(clk), .RN(n4435), .Q(
        \key_mem[8][114] ) );
  DFFRX1 \key_mem_reg[0][113]  ( .D(n1752), .CK(clk), .RN(n4436), .Q(
        \key_mem[0][113] ) );
  DFFRX1 \key_mem_reg[4][113]  ( .D(n2264), .CK(clk), .RN(n4437), .Q(
        \key_mem[4][113] ) );
  DFFRX1 \key_mem_reg[8][113]  ( .D(n2776), .CK(clk), .RN(n4437), .Q(
        \key_mem[8][113] ) );
  DFFRX1 \key_mem_reg[0][112]  ( .D(n1753), .CK(clk), .RN(n4438), .Q(
        \key_mem[0][112] ) );
  DFFRX1 \key_mem_reg[4][112]  ( .D(n2265), .CK(clk), .RN(n4438), .Q(
        \key_mem[4][112] ) );
  DFFRX1 \key_mem_reg[8][112]  ( .D(n2777), .CK(clk), .RN(n4439), .Q(
        \key_mem[8][112] ) );
  DFFRX1 \key_mem_reg[0][111]  ( .D(n1754), .CK(clk), .RN(n4440), .Q(
        \key_mem[0][111] ) );
  DFFRX1 \key_mem_reg[4][111]  ( .D(n2266), .CK(clk), .RN(n4440), .Q(
        \key_mem[4][111] ) );
  DFFRX1 \key_mem_reg[8][111]  ( .D(n2778), .CK(clk), .RN(n4417), .Q(
        \key_mem[8][111] ) );
  DFFRX1 \key_mem_reg[0][110]  ( .D(n1755), .CK(clk), .RN(n4418), .Q(
        \key_mem[0][110] ) );
  DFFRX1 \key_mem_reg[4][110]  ( .D(n2267), .CK(clk), .RN(n4438), .Q(
        \key_mem[4][110] ) );
  DFFRX1 \key_mem_reg[8][110]  ( .D(n2779), .CK(clk), .RN(n4435), .Q(
        \key_mem[8][110] ) );
  DFFRX1 \key_mem_reg[0][109]  ( .D(n1756), .CK(clk), .RN(n4419), .Q(
        \key_mem[0][109] ) );
  DFFRX1 \key_mem_reg[4][109]  ( .D(n2268), .CK(clk), .RN(n4419), .Q(
        \key_mem[4][109] ) );
  DFFRX1 \key_mem_reg[8][109]  ( .D(n2780), .CK(clk), .RN(n4420), .Q(
        \key_mem[8][109] ) );
  DFFRX1 \key_mem_reg[0][108]  ( .D(n1757), .CK(clk), .RN(n4421), .Q(
        \key_mem[0][108] ) );
  DFFRX1 \key_mem_reg[4][108]  ( .D(n2269), .CK(clk), .RN(n4421), .Q(
        \key_mem[4][108] ) );
  DFFRX1 \key_mem_reg[8][108]  ( .D(n2781), .CK(clk), .RN(n4422), .Q(
        \key_mem[8][108] ) );
  DFFRX1 \key_mem_reg[0][107]  ( .D(n1758), .CK(clk), .RN(n4465), .Q(
        \key_mem[0][107] ) );
  DFFRX1 \key_mem_reg[4][107]  ( .D(n2270), .CK(clk), .RN(n4462), .Q(
        \key_mem[4][107] ) );
  DFFRX1 \key_mem_reg[8][107]  ( .D(n2782), .CK(clk), .RN(n4463), .Q(
        \key_mem[8][107] ) );
  DFFRX1 \key_mem_reg[0][106]  ( .D(n1759), .CK(clk), .RN(n4473), .Q(
        \key_mem[0][106] ) );
  DFFRX1 \key_mem_reg[4][106]  ( .D(n2271), .CK(clk), .RN(n4423), .Q(
        \key_mem[4][106] ) );
  DFFRX1 \key_mem_reg[8][106]  ( .D(n2783), .CK(clk), .RN(n4423), .Q(
        \key_mem[8][106] ) );
  DFFRX1 \key_mem_reg[0][105]  ( .D(n1760), .CK(clk), .RN(n4424), .Q(
        \key_mem[0][105] ) );
  DFFRX1 \key_mem_reg[4][105]  ( .D(n2272), .CK(clk), .RN(n4425), .Q(
        \key_mem[4][105] ) );
  DFFRX1 \key_mem_reg[8][105]  ( .D(n2784), .CK(clk), .RN(n4425), .Q(
        \key_mem[8][105] ) );
  DFFRX1 \key_mem_reg[0][104]  ( .D(n1761), .CK(clk), .RN(n4426), .Q(
        \key_mem[0][104] ) );
  DFFRX1 \key_mem_reg[4][104]  ( .D(n2273), .CK(clk), .RN(n4426), .Q(
        \key_mem[4][104] ) );
  DFFRX1 \key_mem_reg[8][104]  ( .D(n2785), .CK(clk), .RN(n4427), .Q(
        \key_mem[8][104] ) );
  DFFRX1 \key_mem_reg[0][103]  ( .D(n1762), .CK(clk), .RN(n4428), .Q(
        \key_mem[0][103] ) );
  DFFRX1 \key_mem_reg[4][103]  ( .D(n2274), .CK(clk), .RN(n4428), .Q(
        \key_mem[4][103] ) );
  DFFRX1 \key_mem_reg[8][103]  ( .D(n2786), .CK(clk), .RN(n4429), .Q(
        \key_mem[8][103] ) );
  DFFRX1 \key_mem_reg[0][102]  ( .D(n1763), .CK(clk), .RN(n4456), .Q(
        \key_mem[0][102] ) );
  DFFRX1 \key_mem_reg[4][102]  ( .D(n2275), .CK(clk), .RN(n4456), .Q(
        \key_mem[4][102] ) );
  DFFRX1 \key_mem_reg[8][102]  ( .D(n2787), .CK(clk), .RN(n4456), .Q(
        \key_mem[8][102] ) );
  DFFRX1 \key_mem_reg[0][101]  ( .D(n1764), .CK(clk), .RN(n4457), .Q(
        \key_mem[0][101] ) );
  DFFRX1 \key_mem_reg[4][101]  ( .D(n2276), .CK(clk), .RN(n4458), .Q(
        \key_mem[4][101] ) );
  DFFRX1 \key_mem_reg[8][101]  ( .D(n2788), .CK(clk), .RN(n4458), .Q(
        \key_mem[8][101] ) );
  DFFRX1 \key_mem_reg[0][100]  ( .D(n1765), .CK(clk), .RN(n4459), .Q(
        \key_mem[0][100] ) );
  DFFRX1 \key_mem_reg[4][100]  ( .D(n2277), .CK(clk), .RN(n4459), .Q(
        \key_mem[4][100] ) );
  DFFRX1 \key_mem_reg[8][100]  ( .D(n2789), .CK(clk), .RN(n4460), .Q(
        \key_mem[8][100] ) );
  DFFRX1 \key_mem_reg[0][99]  ( .D(n1766), .CK(clk), .RN(n4473), .Q(
        \key_mem[0][99] ) );
  DFFRX1 \key_mem_reg[4][99]  ( .D(n2278), .CK(clk), .RN(n4472), .Q(
        \key_mem[4][99] ) );
  DFFRX1 \key_mem_reg[8][99]  ( .D(n2790), .CK(clk), .RN(n4461), .Q(
        \key_mem[8][99] ) );
  DFFRX1 \key_mem_reg[0][98]  ( .D(n1767), .CK(clk), .RN(n4462), .Q(
        \key_mem[0][98] ) );
  DFFRX1 \key_mem_reg[4][98]  ( .D(n2279), .CK(clk), .RN(n4462), .Q(
        \key_mem[4][98] ) );
  DFFRX1 \key_mem_reg[8][98]  ( .D(n2791), .CK(clk), .RN(n4463), .Q(
        \key_mem[8][98] ) );
  DFFRX1 \key_mem_reg[0][97]  ( .D(n1768), .CK(clk), .RN(n4463), .Q(
        \key_mem[0][97] ) );
  DFFRX1 \key_mem_reg[4][97]  ( .D(n2280), .CK(clk), .RN(n4464), .Q(
        \key_mem[4][97] ) );
  DFFRX1 \key_mem_reg[8][97]  ( .D(n2792), .CK(clk), .RN(n4464), .Q(
        \key_mem[8][97] ) );
  DFFRX1 \key_mem_reg[0][96]  ( .D(n1769), .CK(clk), .RN(n4465), .Q(
        \key_mem[0][96] ) );
  DFFRX1 \key_mem_reg[4][96]  ( .D(n2281), .CK(clk), .RN(n4466), .Q(
        \key_mem[4][96] ) );
  DFFRX1 \key_mem_reg[8][96]  ( .D(n2793), .CK(clk), .RN(n4466), .Q(
        \key_mem[8][96] ) );
  DFFRX1 \key_mem_reg[0][87]  ( .D(n1778), .CK(clk), .RN(n4467), .Q(
        \key_mem[0][87] ) );
  DFFRX1 \key_mem_reg[4][87]  ( .D(n2290), .CK(clk), .RN(n4467), .Q(
        \key_mem[4][87] ) );
  DFFRX1 \key_mem_reg[8][87]  ( .D(n2802), .CK(clk), .RN(n4468), .Q(
        \key_mem[8][87] ) );
  DFFRX1 \key_mem_reg[0][86]  ( .D(n1779), .CK(clk), .RN(n4469), .Q(
        \key_mem[0][86] ) );
  DFFRX1 \key_mem_reg[4][86]  ( .D(n2291), .CK(clk), .RN(n4469), .Q(
        \key_mem[4][86] ) );
  DFFRX1 \key_mem_reg[8][86]  ( .D(n2803), .CK(clk), .RN(n4448), .Q(
        \key_mem[8][86] ) );
  DFFRX1 \key_mem_reg[0][85]  ( .D(n1780), .CK(clk), .RN(n4441), .Q(
        \key_mem[0][85] ) );
  DFFRX1 \key_mem_reg[4][85]  ( .D(n2292), .CK(clk), .RN(n4442), .Q(
        \key_mem[4][85] ) );
  DFFRX1 \key_mem_reg[8][85]  ( .D(n2804), .CK(clk), .RN(n4442), .Q(
        \key_mem[8][85] ) );
  DFFRX1 \key_mem_reg[0][84]  ( .D(n1781), .CK(clk), .RN(n4443), .Q(
        \key_mem[0][84] ) );
  DFFRX1 \key_mem_reg[4][84]  ( .D(n2293), .CK(clk), .RN(n4443), .Q(
        \key_mem[4][84] ) );
  DFFRX1 \key_mem_reg[8][84]  ( .D(n2805), .CK(clk), .RN(n4444), .Q(
        \key_mem[8][84] ) );
  DFFRX1 \key_mem_reg[0][83]  ( .D(n1782), .CK(clk), .RN(n4445), .Q(
        \key_mem[0][83] ) );
  DFFRX1 \key_mem_reg[4][83]  ( .D(n2294), .CK(clk), .RN(n4445), .Q(
        \key_mem[4][83] ) );
  DFFRX1 \key_mem_reg[8][83]  ( .D(n2806), .CK(clk), .RN(n4446), .Q(
        \key_mem[8][83] ) );
  DFFRX1 \key_mem_reg[0][82]  ( .D(n1783), .CK(clk), .RN(n4446), .Q(
        \key_mem[0][82] ) );
  DFFRX1 \key_mem_reg[4][82]  ( .D(n2295), .CK(clk), .RN(n4447), .Q(
        \key_mem[4][82] ) );
  DFFRX1 \key_mem_reg[8][82]  ( .D(n2807), .CK(clk), .RN(n4447), .Q(
        \key_mem[8][82] ) );
  DFFRX1 \key_mem_reg[0][81]  ( .D(n1784), .CK(clk), .RN(n4448), .Q(
        \key_mem[0][81] ) );
  DFFRX1 \key_mem_reg[4][81]  ( .D(n2296), .CK(clk), .RN(n4449), .Q(
        \key_mem[4][81] ) );
  DFFRX1 \key_mem_reg[8][81]  ( .D(n2808), .CK(clk), .RN(n4449), .Q(
        \key_mem[8][81] ) );
  DFFRX1 \key_mem_reg[0][80]  ( .D(n1785), .CK(clk), .RN(n4450), .Q(
        \key_mem[0][80] ) );
  DFFRX1 \key_mem_reg[4][80]  ( .D(n2297), .CK(clk), .RN(n4450), .Q(
        \key_mem[4][80] ) );
  DFFRX1 \key_mem_reg[8][80]  ( .D(n2809), .CK(clk), .RN(n4451), .Q(
        \key_mem[8][80] ) );
  DFFRX1 \key_mem_reg[0][79]  ( .D(n1786), .CK(clk), .RN(n4452), .Q(
        \key_mem[0][79] ) );
  DFFRX1 \key_mem_reg[4][79]  ( .D(n2298), .CK(clk), .RN(n4452), .Q(
        \key_mem[4][79] ) );
  DFFRX1 \key_mem_reg[8][79]  ( .D(n2810), .CK(clk), .RN(n4453), .Q(
        \key_mem[8][79] ) );
  DFFRX1 \key_mem_reg[0][78]  ( .D(n1787), .CK(clk), .RN(n4454), .Q(
        \key_mem[0][78] ) );
  DFFRX1 \key_mem_reg[4][78]  ( .D(n2299), .CK(clk), .RN(n4454), .Q(
        \key_mem[4][78] ) );
  DFFRX1 \key_mem_reg[8][78]  ( .D(n2811), .CK(clk), .RN(n4454), .Q(
        \key_mem[8][78] ) );
  DFFRX1 \key_mem_reg[0][77]  ( .D(n1788), .CK(clk), .RN(n4455), .Q(
        \key_mem[0][77] ) );
  DFFRX1 \key_mem_reg[4][77]  ( .D(n2300), .CK(clk), .RN(n4380), .Q(
        \key_mem[4][77] ) );
  DFFRX1 \key_mem_reg[8][77]  ( .D(n2812), .CK(clk), .RN(n4373), .Q(
        \key_mem[8][77] ) );
  DFFRX1 \key_mem_reg[0][76]  ( .D(n1789), .CK(clk), .RN(n4374), .Q(
        \key_mem[0][76] ) );
  DFFRX1 \key_mem_reg[4][76]  ( .D(n2301), .CK(clk), .RN(n4374), .Q(
        \key_mem[4][76] ) );
  DFFRX1 \key_mem_reg[8][76]  ( .D(n2813), .CK(clk), .RN(n4375), .Q(
        \key_mem[8][76] ) );
  DFFRX1 \key_mem_reg[0][75]  ( .D(n1790), .CK(clk), .RN(n4376), .Q(
        \key_mem[0][75] ) );
  DFFRX1 \key_mem_reg[4][75]  ( .D(n2302), .CK(clk), .RN(n4376), .Q(
        \key_mem[4][75] ) );
  DFFRX1 \key_mem_reg[8][75]  ( .D(n2814), .CK(clk), .RN(n4377), .Q(
        \key_mem[8][75] ) );
  DFFRX1 \key_mem_reg[0][74]  ( .D(n1791), .CK(clk), .RN(n4378), .Q(
        \key_mem[0][74] ) );
  DFFRX1 \key_mem_reg[4][74]  ( .D(n2303), .CK(clk), .RN(n4378), .Q(
        \key_mem[4][74] ) );
  DFFRX1 \key_mem_reg[8][74]  ( .D(n2815), .CK(clk), .RN(n4378), .Q(
        \key_mem[8][74] ) );
  DFFRX1 \key_mem_reg[0][73]  ( .D(n1792), .CK(clk), .RN(n4379), .Q(
        \key_mem[0][73] ) );
  DFFRX1 \key_mem_reg[4][73]  ( .D(n2304), .CK(clk), .RN(n4380), .Q(
        \key_mem[4][73] ) );
  DFFRX1 \key_mem_reg[8][73]  ( .D(n2816), .CK(clk), .RN(n4380), .Q(
        \key_mem[8][73] ) );
  DFFRX1 \key_mem_reg[0][72]  ( .D(n1793), .CK(clk), .RN(n4381), .Q(
        \key_mem[0][72] ) );
  DFFRX1 \key_mem_reg[4][72]  ( .D(n2305), .CK(clk), .RN(n4382), .Q(
        \key_mem[4][72] ) );
  DFFRX1 \key_mem_reg[8][72]  ( .D(n2817), .CK(clk), .RN(n4382), .Q(
        \key_mem[8][72] ) );
  DFFRX1 \key_mem_reg[0][71]  ( .D(n1794), .CK(clk), .RN(n4383), .Q(
        \key_mem[0][71] ) );
  DFFRX1 \key_mem_reg[4][71]  ( .D(n2306), .CK(clk), .RN(n4383), .Q(
        \key_mem[4][71] ) );
  DFFRX1 \key_mem_reg[8][71]  ( .D(n2818), .CK(clk), .RN(n4384), .Q(
        \key_mem[8][71] ) );
  DFFRX1 \key_mem_reg[0][70]  ( .D(n1795), .CK(clk), .RN(n4385), .Q(
        \key_mem[0][70] ) );
  DFFRX1 \key_mem_reg[4][70]  ( .D(n2307), .CK(clk), .RN(n4385), .Q(
        \key_mem[4][70] ) );
  DFFRX1 \key_mem_reg[8][70]  ( .D(n2819), .CK(clk), .RN(n4386), .Q(
        \key_mem[8][70] ) );
  DFFRX1 \key_mem_reg[0][69]  ( .D(n1796), .CK(clk), .RN(n4386), .Q(
        \key_mem[0][69] ) );
  DFFRX1 \key_mem_reg[4][69]  ( .D(n2308), .CK(clk), .RN(n4387), .Q(
        \key_mem[4][69] ) );
  DFFRX1 \key_mem_reg[8][69]  ( .D(n2820), .CK(clk), .RN(n4387), .Q(
        \key_mem[8][69] ) );
  DFFRX1 \key_mem_reg[0][68]  ( .D(n1797), .CK(clk), .RN(n4504), .Q(
        \key_mem[0][68] ) );
  DFFRX1 \key_mem_reg[4][68]  ( .D(n2309), .CK(clk), .RN(n4503), .Q(
        \key_mem[4][68] ) );
  DFFRX1 \key_mem_reg[8][68]  ( .D(n2821), .CK(clk), .RN(n4383), .Q(
        \key_mem[8][68] ) );
  DFFRX1 \key_mem_reg[0][67]  ( .D(n1798), .CK(clk), .RN(n4388), .Q(
        \key_mem[0][67] ) );
  DFFRX1 \key_mem_reg[4][67]  ( .D(n2310), .CK(clk), .RN(n4387), .Q(
        \key_mem[4][67] ) );
  DFFRX1 \key_mem_reg[8][67]  ( .D(n2822), .CK(clk), .RN(n4377), .Q(
        \key_mem[8][67] ) );
  DFFRX1 \key_mem_reg[0][66]  ( .D(n1799), .CK(clk), .RN(n4406), .Q(
        \key_mem[0][66] ) );
  DFFRX1 \key_mem_reg[4][66]  ( .D(n2311), .CK(clk), .RN(n4405), .Q(
        \key_mem[4][66] ) );
  DFFRX1 \key_mem_reg[8][66]  ( .D(n2823), .CK(clk), .RN(n4404), .Q(
        \key_mem[8][66] ) );
  DFFRX1 \key_mem_reg[0][65]  ( .D(n1800), .CK(clk), .RN(n4397), .Q(
        \key_mem[0][65] ) );
  DFFRX1 \key_mem_reg[4][65]  ( .D(n2312), .CK(clk), .RN(n4453), .Q(
        \key_mem[4][65] ) );
  DFFRX1 \key_mem_reg[8][65]  ( .D(n2824), .CK(clk), .RN(n4454), .Q(
        \key_mem[8][65] ) );
  DFFRX1 \key_mem_reg[0][64]  ( .D(n1801), .CK(clk), .RN(n4445), .Q(
        \key_mem[0][64] ) );
  DFFRX1 \key_mem_reg[4][64]  ( .D(n2313), .CK(clk), .RN(n4420), .Q(
        \key_mem[4][64] ) );
  DFFRX1 \key_mem_reg[8][64]  ( .D(n2825), .CK(clk), .RN(n4418), .Q(
        \key_mem[8][64] ) );
  DFFRX1 \key_mem_reg[0][55]  ( .D(n1810), .CK(clk), .RN(n4499), .Q(
        \key_mem[0][55] ) );
  DFFRX1 \key_mem_reg[4][55]  ( .D(n2322), .CK(clk), .RN(n4526), .Q(
        \key_mem[4][55] ) );
  DFFRX1 \key_mem_reg[8][55]  ( .D(n2834), .CK(clk), .RN(n4553), .Q(
        \key_mem[8][55] ) );
  DFFRX1 \key_mem_reg[0][54]  ( .D(n1811), .CK(clk), .RN(n4540), .Q(
        \key_mem[0][54] ) );
  DFFRX1 \key_mem_reg[4][54]  ( .D(n2323), .CK(clk), .RN(n4539), .Q(
        \key_mem[4][54] ) );
  DFFRX1 \key_mem_reg[8][54]  ( .D(n2835), .CK(clk), .RN(n4370), .Q(
        \key_mem[8][54] ) );
  DFFRX1 \key_mem_reg[0][53]  ( .D(n1812), .CK(clk), .RN(n4370), .Q(
        \key_mem[0][53] ) );
  DFFRX1 \key_mem_reg[4][53]  ( .D(n2324), .CK(clk), .RN(n4371), .Q(
        \key_mem[4][53] ) );
  DFFRX1 \key_mem_reg[8][53]  ( .D(n2836), .CK(clk), .RN(n4371), .Q(
        \key_mem[8][53] ) );
  DFFRX1 \key_mem_reg[0][52]  ( .D(n1813), .CK(clk), .RN(n4372), .Q(
        \key_mem[0][52] ) );
  DFFRX1 \key_mem_reg[4][52]  ( .D(n2325), .CK(clk), .RN(n4373), .Q(
        \key_mem[4][52] ) );
  DFFRX1 \key_mem_reg[8][52]  ( .D(n2837), .CK(clk), .RN(n4403), .Q(
        \key_mem[8][52] ) );
  DFFRX1 \key_mem_reg[0][51]  ( .D(n1814), .CK(clk), .RN(n4404), .Q(
        \key_mem[0][51] ) );
  DFFRX1 \key_mem_reg[4][51]  ( .D(n2326), .CK(clk), .RN(n4404), .Q(
        \key_mem[4][51] ) );
  DFFRX1 \key_mem_reg[8][51]  ( .D(n2838), .CK(clk), .RN(n4405), .Q(
        \key_mem[8][51] ) );
  DFFRX1 \key_mem_reg[0][50]  ( .D(n1815), .CK(clk), .RN(n4406), .Q(
        \key_mem[0][50] ) );
  DFFRX1 \key_mem_reg[4][50]  ( .D(n2327), .CK(clk), .RN(n4406), .Q(
        \key_mem[4][50] ) );
  DFFRX1 \key_mem_reg[8][50]  ( .D(n2839), .CK(clk), .RN(n4407), .Q(
        \key_mem[8][50] ) );
  DFFRX1 \key_mem_reg[0][49]  ( .D(n1816), .CK(clk), .RN(n4408), .Q(
        \key_mem[0][49] ) );
  DFFRX1 \key_mem_reg[4][49]  ( .D(n2328), .CK(clk), .RN(n4408), .Q(
        \key_mem[4][49] ) );
  DFFRX1 \key_mem_reg[8][49]  ( .D(n2840), .CK(clk), .RN(n4408), .Q(
        \key_mem[8][49] ) );
  DFFRX1 \key_mem_reg[0][47]  ( .D(n1818), .CK(clk), .RN(n4411), .Q(
        \key_mem[0][47] ) );
  DFFRX1 \key_mem_reg[4][47]  ( .D(n2330), .CK(clk), .RN(n4412), .Q(
        \key_mem[4][47] ) );
  DFFRX1 \key_mem_reg[8][47]  ( .D(n2842), .CK(clk), .RN(n4412), .Q(
        \key_mem[8][47] ) );
  DFFRX1 \key_mem_reg[0][46]  ( .D(n1819), .CK(clk), .RN(n4413), .Q(
        \key_mem[0][46] ) );
  DFFRX1 \key_mem_reg[4][46]  ( .D(n2331), .CK(clk), .RN(n4413), .Q(
        \key_mem[4][46] ) );
  DFFRX1 \key_mem_reg[8][46]  ( .D(n2843), .CK(clk), .RN(n4409), .Q(
        \key_mem[8][46] ) );
  DFFRX1 \key_mem_reg[0][45]  ( .D(n1820), .CK(clk), .RN(n4414), .Q(
        \key_mem[0][45] ) );
  DFFRX1 \key_mem_reg[4][45]  ( .D(n2332), .CK(clk), .RN(n4414), .Q(
        \key_mem[4][45] ) );
  DFFRX1 \key_mem_reg[8][45]  ( .D(n2844), .CK(clk), .RN(n4415), .Q(
        \key_mem[8][45] ) );
  DFFRX1 \key_mem_reg[0][44]  ( .D(n1821), .CK(clk), .RN(n4415), .Q(
        \key_mem[0][44] ) );
  DFFRX1 \key_mem_reg[4][44]  ( .D(n2333), .CK(clk), .RN(n4416), .Q(
        \key_mem[4][44] ) );
  DFFRX1 \key_mem_reg[8][44]  ( .D(n2845), .CK(clk), .RN(n4416), .Q(
        \key_mem[8][44] ) );
  DFFRX1 \key_mem_reg[0][43]  ( .D(n1822), .CK(clk), .RN(n4388), .Q(
        \key_mem[0][43] ) );
  DFFRX1 \key_mem_reg[4][43]  ( .D(n2334), .CK(clk), .RN(n4388), .Q(
        \key_mem[4][43] ) );
  DFFRX1 \key_mem_reg[8][43]  ( .D(n2846), .CK(clk), .RN(n4389), .Q(
        \key_mem[8][43] ) );
  DFFRX1 \key_mem_reg[0][42]  ( .D(n1823), .CK(clk), .RN(n4390), .Q(
        \key_mem[0][42] ) );
  DFFRX1 \key_mem_reg[4][42]  ( .D(n2335), .CK(clk), .RN(n4390), .Q(
        \key_mem[4][42] ) );
  DFFRX1 \key_mem_reg[8][42]  ( .D(n2847), .CK(clk), .RN(n4391), .Q(
        \key_mem[8][42] ) );
  DFFRX1 \key_mem_reg[0][41]  ( .D(n1824), .CK(clk), .RN(n4391), .Q(
        \key_mem[0][41] ) );
  DFFRX1 \key_mem_reg[4][41]  ( .D(n2336), .CK(clk), .RN(n4392), .Q(
        \key_mem[4][41] ) );
  DFFRX1 \key_mem_reg[8][41]  ( .D(n2848), .CK(clk), .RN(n4392), .Q(
        \key_mem[8][41] ) );
  DFFRX1 \key_mem_reg[0][40]  ( .D(n1825), .CK(clk), .RN(n4393), .Q(
        \key_mem[0][40] ) );
  DFFRX1 \key_mem_reg[4][40]  ( .D(n2337), .CK(clk), .RN(n4394), .Q(
        \key_mem[4][40] ) );
  DFFRX1 \key_mem_reg[8][40]  ( .D(n2849), .CK(clk), .RN(n4394), .Q(
        \key_mem[8][40] ) );
  DFFRX1 \key_mem_reg[0][39]  ( .D(n1826), .CK(clk), .RN(n4395), .Q(
        \key_mem[0][39] ) );
  DFFRX1 \key_mem_reg[4][39]  ( .D(n2338), .CK(clk), .RN(n4395), .Q(
        \key_mem[4][39] ) );
  DFFRX1 \key_mem_reg[8][39]  ( .D(n2850), .CK(clk), .RN(n4396), .Q(
        \key_mem[8][39] ) );
  DFFRX1 \key_mem_reg[0][38]  ( .D(n1827), .CK(clk), .RN(n4397), .Q(
        \key_mem[0][38] ) );
  DFFRX1 \key_mem_reg[4][38]  ( .D(n2339), .CK(clk), .RN(n4397), .Q(
        \key_mem[4][38] ) );
  DFFRX1 \key_mem_reg[8][38]  ( .D(n2851), .CK(clk), .RN(n4398), .Q(
        \key_mem[8][38] ) );
  DFFRX1 \key_mem_reg[0][37]  ( .D(n1828), .CK(clk), .RN(n4399), .Q(
        \key_mem[0][37] ) );
  DFFRX1 \key_mem_reg[4][37]  ( .D(n2340), .CK(clk), .RN(n4399), .Q(
        \key_mem[4][37] ) );
  DFFRX1 \key_mem_reg[8][37]  ( .D(n2852), .CK(clk), .RN(n4399), .Q(
        \key_mem[8][37] ) );
  DFFRX1 \key_mem_reg[0][36]  ( .D(n1829), .CK(clk), .RN(n4400), .Q(
        \key_mem[0][36] ) );
  DFFRX1 \key_mem_reg[4][36]  ( .D(n2341), .CK(clk), .RN(n4401), .Q(
        \key_mem[4][36] ) );
  DFFRX1 \key_mem_reg[8][36]  ( .D(n2853), .CK(clk), .RN(n4401), .Q(
        \key_mem[8][36] ) );
  DFFRX1 \key_mem_reg[0][35]  ( .D(n1830), .CK(clk), .RN(n4402), .Q(
        \key_mem[0][35] ) );
  DFFRX1 \key_mem_reg[4][35]  ( .D(n2342), .CK(clk), .RN(n4402), .Q(
        \key_mem[4][35] ) );
  DFFRX1 \key_mem_reg[8][35]  ( .D(n2854), .CK(clk), .RN(n4403), .Q(
        \key_mem[8][35] ) );
  DFFRX1 \key_mem_reg[0][34]  ( .D(n1831), .CK(clk), .RN(n4542), .Q(
        \key_mem[0][34] ) );
  DFFRX1 \key_mem_reg[4][34]  ( .D(n2343), .CK(clk), .RN(n4542), .Q(
        \key_mem[4][34] ) );
  DFFRX1 \key_mem_reg[8][34]  ( .D(n2855), .CK(clk), .RN(n4543), .Q(
        \key_mem[8][34] ) );
  DFFRX1 \key_mem_reg[0][33]  ( .D(n1832), .CK(clk), .RN(n4543), .Q(
        \key_mem[0][33] ) );
  DFFRX1 \key_mem_reg[4][33]  ( .D(n2344), .CK(clk), .RN(n4544), .Q(
        \key_mem[4][33] ) );
  DFFRX1 \key_mem_reg[8][33]  ( .D(n2856), .CK(clk), .RN(n4544), .Q(
        \key_mem[8][33] ) );
  DFFRX1 \key_mem_reg[0][32]  ( .D(n1833), .CK(clk), .RN(n4545), .Q(
        \key_mem[0][32] ) );
  DFFRX1 \key_mem_reg[4][32]  ( .D(n2345), .CK(clk), .RN(n4546), .Q(
        \key_mem[4][32] ) );
  DFFRX1 \key_mem_reg[8][32]  ( .D(n2857), .CK(clk), .RN(n4546), .Q(
        \key_mem[8][32] ) );
  DFFRX1 \key_mem_reg[0][23]  ( .D(n1842), .CK(clk), .RN(n4547), .Q(
        \key_mem[0][23] ) );
  DFFRX1 \key_mem_reg[4][23]  ( .D(n2354), .CK(clk), .RN(n4547), .Q(
        \key_mem[4][23] ) );
  DFFRX1 \key_mem_reg[8][23]  ( .D(n2866), .CK(clk), .RN(n4548), .Q(
        \key_mem[8][23] ) );
  DFFRX1 \key_mem_reg[0][22]  ( .D(n1843), .CK(clk), .RN(n4549), .Q(
        \key_mem[0][22] ) );
  DFFRX1 \key_mem_reg[4][22]  ( .D(n2355), .CK(clk), .RN(n4549), .Q(
        \key_mem[4][22] ) );
  DFFRX1 \key_mem_reg[8][22]  ( .D(n2867), .CK(clk), .RN(n4550), .Q(
        \key_mem[8][22] ) );
  DFFRX1 \key_mem_reg[0][21]  ( .D(n1844), .CK(clk), .RN(n4551), .Q(
        \key_mem[0][21] ) );
  DFFRX1 \key_mem_reg[4][21]  ( .D(n2356), .CK(clk), .RN(n4551), .Q(
        \key_mem[4][21] ) );
  DFFRX1 \key_mem_reg[8][21]  ( .D(n2868), .CK(clk), .RN(n4551), .Q(
        \key_mem[8][21] ) );
  DFFRX1 \key_mem_reg[0][20]  ( .D(n1845), .CK(clk), .RN(n4552), .Q(
        \key_mem[0][20] ) );
  DFFRX1 \key_mem_reg[4][20]  ( .D(n2357), .CK(clk), .RN(n4553), .Q(
        \key_mem[4][20] ) );
  DFFRX1 \key_mem_reg[8][20]  ( .D(n2869), .CK(clk), .RN(n4553), .Q(
        \key_mem[8][20] ) );
  DFFRX1 \key_mem_reg[0][19]  ( .D(n1846), .CK(clk), .RN(n4421), .Q(
        \key_mem[0][19] ) );
  DFFRX1 \key_mem_reg[4][19]  ( .D(n2358), .CK(clk), .RN(n4422), .Q(
        \key_mem[4][19] ) );
  DFFRX1 \key_mem_reg[8][19]  ( .D(n2870), .CK(clk), .RN(n4480), .Q(
        \key_mem[8][19] ) );
  DFFRX1 \key_mem_reg[0][18]  ( .D(n1847), .CK(clk), .RN(n4554), .Q(
        \key_mem[0][18] ) );
  DFFRX1 \key_mem_reg[4][18]  ( .D(n2359), .CK(clk), .RN(n4554), .Q(
        \key_mem[4][18] ) );
  DFFRX1 \key_mem_reg[8][18]  ( .D(n2871), .CK(clk), .RN(n4526), .Q(
        \key_mem[8][18] ) );
  DFFRX1 \key_mem_reg[0][17]  ( .D(n1848), .CK(clk), .RN(n4527), .Q(
        \key_mem[0][17] ) );
  DFFRX1 \key_mem_reg[4][17]  ( .D(n2360), .CK(clk), .RN(n4528), .Q(
        \key_mem[4][17] ) );
  DFFRX1 \key_mem_reg[8][17]  ( .D(n2872), .CK(clk), .RN(n4528), .Q(
        \key_mem[8][17] ) );
  DFFRX1 \key_mem_reg[0][16]  ( .D(n1849), .CK(clk), .RN(n4529), .Q(
        \key_mem[0][16] ) );
  DFFRX1 \key_mem_reg[4][16]  ( .D(n2361), .CK(clk), .RN(n4529), .Q(
        \key_mem[4][16] ) );
  DFFRX1 \key_mem_reg[8][16]  ( .D(n2873), .CK(clk), .RN(n4530), .Q(
        \key_mem[8][16] ) );
  DFFRX1 \key_mem_reg[0][15]  ( .D(n1850), .CK(clk), .RN(n4531), .Q(
        \key_mem[0][15] ) );
  DFFRX1 \key_mem_reg[4][15]  ( .D(n2362), .CK(clk), .RN(n4531), .Q(
        \key_mem[4][15] ) );
  DFFRX1 \key_mem_reg[8][15]  ( .D(n2874), .CK(clk), .RN(n4532), .Q(
        \key_mem[8][15] ) );
  DFFRX1 \key_mem_reg[0][14]  ( .D(n1851), .CK(clk), .RN(n4533), .Q(
        \key_mem[0][14] ) );
  DFFRX1 \key_mem_reg[4][14]  ( .D(n2363), .CK(clk), .RN(n4533), .Q(
        \key_mem[4][14] ) );
  DFFRX1 \key_mem_reg[8][14]  ( .D(n2875), .CK(clk), .RN(n4533), .Q(
        \key_mem[8][14] ) );
  DFFRX1 \key_mem_reg[0][13]  ( .D(n1852), .CK(clk), .RN(n4534), .Q(
        \key_mem[0][13] ) );
  DFFRX1 \key_mem_reg[4][13]  ( .D(n2364), .CK(clk), .RN(n4535), .Q(
        \key_mem[4][13] ) );
  DFFRX1 \key_mem_reg[8][13]  ( .D(n2876), .CK(clk), .RN(n4535), .Q(
        \key_mem[8][13] ) );
  DFFRX1 \key_mem_reg[0][12]  ( .D(n1853), .CK(clk), .RN(n4536), .Q(
        \key_mem[0][12] ) );
  DFFRX1 \key_mem_reg[4][12]  ( .D(n2365), .CK(clk), .RN(n4537), .Q(
        \key_mem[4][12] ) );
  DFFRX1 \key_mem_reg[8][12]  ( .D(n2877), .CK(clk), .RN(n4537), .Q(
        \key_mem[8][12] ) );
  DFFRX1 \key_mem_reg[0][11]  ( .D(n1854), .CK(clk), .RN(n4538), .Q(
        \key_mem[0][11] ) );
  DFFRX1 \key_mem_reg[4][11]  ( .D(n2366), .CK(clk), .RN(n4538), .Q(
        \key_mem[4][11] ) );
  DFFRX1 \key_mem_reg[8][11]  ( .D(n2878), .CK(clk), .RN(n4539), .Q(
        \key_mem[8][11] ) );
  DFFRX1 \key_mem_reg[0][10]  ( .D(n1855), .CK(clk), .RN(n4540), .Q(
        \key_mem[0][10] ) );
  DFFRX1 \key_mem_reg[4][10]  ( .D(n2367), .CK(clk), .RN(n4540), .Q(
        \key_mem[4][10] ) );
  DFFRX1 \key_mem_reg[8][10]  ( .D(n2879), .CK(clk), .RN(n4541), .Q(
        \key_mem[8][10] ) );
  DFFRX1 \key_mem_reg[0][9]  ( .D(n1856), .CK(clk), .RN(n4502), .Q(
        \key_mem[0][9] ) );
  DFFRX1 \key_mem_reg[4][9]  ( .D(n2368), .CK(clk), .RN(n4536), .Q(
        \key_mem[4][9] ) );
  DFFRX1 \key_mem_reg[8][9]  ( .D(n2880), .CK(clk), .RN(n4501), .Q(
        \key_mem[8][9] ) );
  DFFRX1 \key_mem_reg[0][8]  ( .D(n1857), .CK(clk), .RN(n4529), .Q(
        \key_mem[0][8] ) );
  DFFRX1 \key_mem_reg[4][8]  ( .D(n2369), .CK(clk), .RN(n4497), .Q(
        \key_mem[4][8] ) );
  DFFRX1 \key_mem_reg[8][8]  ( .D(n2881), .CK(clk), .RN(n4521), .Q(
        \key_mem[8][8] ) );
  DFFRX1 \key_mem_reg[0][7]  ( .D(n1858), .CK(clk), .RN(n4559), .Q(
        \key_mem[0][7] ) );
  DFFRX1 \key_mem_reg[4][7]  ( .D(n2370), .CK(clk), .RN(n4559), .Q(
        \key_mem[4][7] ) );
  DFFRX1 \key_mem_reg[8][7]  ( .D(n2882), .CK(clk), .RN(n4560), .Q(
        \key_mem[8][7] ) );
  DFFRX1 \key_mem_reg[0][6]  ( .D(n1859), .CK(clk), .RN(n4561), .Q(
        \key_mem[0][6] ) );
  DFFRX1 \key_mem_reg[4][6]  ( .D(n2371), .CK(clk), .RN(n4561), .Q(
        \key_mem[4][6] ) );
  DFFRX1 \key_mem_reg[8][6]  ( .D(n2883), .CK(clk), .RN(n4562), .Q(
        \key_mem[8][6] ) );
  DFFRX1 \key_mem_reg[0][5]  ( .D(n1860), .CK(clk), .RN(n4376), .Q(
        \key_mem[0][5] ) );
  DFFRX1 \key_mem_reg[4][5]  ( .D(n2372), .CK(clk), .RN(n4440), .Q(
        \key_mem[4][5] ) );
  DFFRX1 \key_mem_reg[8][5]  ( .D(n2884), .CK(clk), .RN(n4434), .Q(
        \key_mem[8][5] ) );
  DFFRX1 \key_mem_reg[0][4]  ( .D(n1861), .CK(clk), .RN(n4429), .Q(
        \key_mem[0][4] ) );
  DFFRX1 \key_mem_reg[4][4]  ( .D(n2373), .CK(clk), .RN(n4415), .Q(
        \key_mem[4][4] ) );
  DFFRX1 \key_mem_reg[8][4]  ( .D(n2885), .CK(clk), .RN(n4416), .Q(
        \key_mem[8][4] ) );
  DFFRX1 \key_mem_reg[0][3]  ( .D(n1862), .CK(clk), .RN(n4466), .Q(
        \key_mem[0][3] ) );
  DFFRX1 \key_mem_reg[4][3]  ( .D(n2374), .CK(clk), .RN(n4380), .Q(
        \key_mem[4][3] ) );
  DFFRX1 \key_mem_reg[8][3]  ( .D(n2886), .CK(clk), .RN(n4383), .Q(
        \key_mem[8][3] ) );
  DFFRX1 \key_mem_reg[0][2]  ( .D(n1863), .CK(clk), .RN(n4375), .Q(
        \key_mem[0][2] ) );
  DFFRX1 \key_mem_reg[4][2]  ( .D(n2375), .CK(clk), .RN(n4467), .Q(
        \key_mem[4][2] ) );
  DFFRX1 \key_mem_reg[8][2]  ( .D(n2887), .CK(clk), .RN(n4563), .Q(
        \key_mem[8][2] ) );
  DFFRX1 \key_mem_reg[0][1]  ( .D(n1864), .CK(clk), .RN(n4564), .Q(
        \key_mem[0][1] ) );
  DFFRX1 \key_mem_reg[4][1]  ( .D(n2376), .CK(clk), .RN(n4564), .Q(
        \key_mem[4][1] ) );
  DFFRX1 \key_mem_reg[8][1]  ( .D(n2888), .CK(clk), .RN(n4554), .Q(
        \key_mem[8][1] ) );
  DFFRX1 \key_mem_reg[0][0]  ( .D(n1865), .CK(clk), .RN(n4555), .Q(
        \key_mem[0][0] ) );
  DFFRX1 \key_mem_reg[4][0]  ( .D(n2377), .CK(clk), .RN(n4556), .Q(
        \key_mem[4][0] ) );
  DFFRX1 \key_mem_reg[8][0]  ( .D(n2889), .CK(clk), .RN(n4556), .Q(
        \key_mem[8][0] ) );
  DFFRX1 \key_mem_reg[0][127]  ( .D(n1738), .CK(clk), .RN(n4489), .Q(
        \key_mem[0][127] ) );
  DFFRX1 \key_mem_reg[4][127]  ( .D(n2250), .CK(clk), .RN(n4488), .Q(
        \key_mem[4][127] ) );
  DFFRX1 \key_mem_reg[8][127]  ( .D(n2762), .CK(clk), .RN(n4531), .Q(
        \key_mem[8][127] ) );
  DFFRX1 \key_mem_reg[0][95]  ( .D(n1770), .CK(clk), .RN(n4523), .Q(
        \key_mem[0][95] ) );
  DFFRX1 \key_mem_reg[4][95]  ( .D(n2282), .CK(clk), .RN(n4522), .Q(
        \key_mem[4][95] ) );
  DFFRX1 \key_mem_reg[8][95]  ( .D(n2794), .CK(clk), .RN(n4512), .Q(
        \key_mem[8][95] ) );
  DFFRX1 \key_mem_reg[0][63]  ( .D(n1802), .CK(clk), .RN(n4560), .Q(
        \key_mem[0][63] ) );
  DFFRX1 \key_mem_reg[4][63]  ( .D(n2314), .CK(clk), .RN(n4559), .Q(
        \key_mem[4][63] ) );
  DFFRX1 \key_mem_reg[8][63]  ( .D(n2826), .CK(clk), .RN(n4548), .Q(
        \key_mem[8][63] ) );
  DFFRX1 \key_mem_reg[0][31]  ( .D(n1834), .CK(clk), .RN(n4485), .Q(
        \key_mem[0][31] ) );
  DFFRX1 \key_mem_reg[4][31]  ( .D(n2346), .CK(clk), .RN(n4557), .Q(
        \key_mem[4][31] ) );
  DFFRX1 \key_mem_reg[8][31]  ( .D(n2858), .CK(clk), .RN(n4557), .Q(
        \key_mem[8][31] ) );
  DFFRX1 \key_mem_reg[0][120]  ( .D(n1745), .CK(clk), .RN(n4460), .Q(
        \key_mem[0][120] ) );
  DFFRX1 \key_mem_reg[4][120]  ( .D(n2257), .CK(clk), .RN(n4489), .Q(
        \key_mem[4][120] ) );
  DFFRX1 \key_mem_reg[8][120]  ( .D(n2769), .CK(clk), .RN(n4488), .Q(
        \key_mem[8][120] ) );
  DFFRX1 \key_mem_reg[0][88]  ( .D(n1777), .CK(clk), .RN(n4543), .Q(
        \key_mem[0][88] ) );
  DFFRX1 \key_mem_reg[4][88]  ( .D(n2289), .CK(clk), .RN(n4542), .Q(
        \key_mem[4][88] ) );
  DFFRX1 \key_mem_reg[8][88]  ( .D(n2801), .CK(clk), .RN(n4558), .Q(
        \key_mem[8][88] ) );
  DFFRX1 \key_mem_reg[0][56]  ( .D(n1809), .CK(clk), .RN(n4474), .Q(
        \key_mem[0][56] ) );
  DFFRX1 \key_mem_reg[4][56]  ( .D(n2321), .CK(clk), .RN(n4519), .Q(
        \key_mem[4][56] ) );
  DFFRX1 \key_mem_reg[8][56]  ( .D(n2833), .CK(clk), .RN(n4509), .Q(
        \key_mem[8][56] ) );
  DFFRX1 \key_mem_reg[0][24]  ( .D(n1841), .CK(clk), .RN(n4496), .Q(
        \key_mem[0][24] ) );
  DFFRX1 \key_mem_reg[4][24]  ( .D(n2353), .CK(clk), .RN(n4450), .Q(
        \key_mem[4][24] ) );
  DFFRX1 \key_mem_reg[8][24]  ( .D(n2865), .CK(clk), .RN(n4447), .Q(
        \key_mem[8][24] ) );
  DFFRX1 \key_mem_reg[0][122]  ( .D(n1743), .CK(clk), .RN(n4485), .Q(
        \key_mem[0][122] ) );
  DFFRX1 \key_mem_reg[4][122]  ( .D(n2255), .CK(clk), .RN(n4485), .Q(
        \key_mem[4][122] ) );
  DFFRX1 \key_mem_reg[8][122]  ( .D(n2767), .CK(clk), .RN(n4485), .Q(
        \key_mem[8][122] ) );
  DFFRX1 \key_mem_reg[0][90]  ( .D(n1775), .CK(clk), .RN(n4486), .Q(
        \key_mem[0][90] ) );
  DFFRX1 \key_mem_reg[4][90]  ( .D(n2287), .CK(clk), .RN(n4487), .Q(
        \key_mem[4][90] ) );
  DFFRX1 \key_mem_reg[8][90]  ( .D(n2799), .CK(clk), .RN(n4487), .Q(
        \key_mem[8][90] ) );
  DFFRX1 \key_mem_reg[0][58]  ( .D(n1807), .CK(clk), .RN(n4488), .Q(
        \key_mem[0][58] ) );
  DFFRX1 \key_mem_reg[4][58]  ( .D(n2319), .CK(clk), .RN(n4488), .Q(
        \key_mem[4][58] ) );
  DFFRX1 \key_mem_reg[8][58]  ( .D(n2831), .CK(clk), .RN(n4489), .Q(
        \key_mem[8][58] ) );
  DFFRX1 \key_mem_reg[0][26]  ( .D(n1839), .CK(clk), .RN(n4490), .Q(
        \key_mem[0][26] ) );
  DFFRX1 \key_mem_reg[4][26]  ( .D(n2351), .CK(clk), .RN(n4490), .Q(
        \key_mem[4][26] ) );
  DFFRX1 \key_mem_reg[8][26]  ( .D(n2863), .CK(clk), .RN(n4491), .Q(
        \key_mem[8][26] ) );
  DFFRX1 \key_mem_reg[0][123]  ( .D(n1742), .CK(clk), .RN(n4535), .Q(
        \key_mem[0][123] ) );
  DFFRX1 \key_mem_reg[4][123]  ( .D(n2254), .CK(clk), .RN(n4503), .Q(
        \key_mem[4][123] ) );
  DFFRX1 \key_mem_reg[8][123]  ( .D(n2766), .CK(clk), .RN(n4429), .Q(
        \key_mem[8][123] ) );
  DFFRX1 \key_mem_reg[0][91]  ( .D(n1774), .CK(clk), .RN(n4492), .Q(
        \key_mem[0][91] ) );
  DFFRX1 \key_mem_reg[4][91]  ( .D(n2286), .CK(clk), .RN(n4492), .Q(
        \key_mem[4][91] ) );
  DFFRX1 \key_mem_reg[8][91]  ( .D(n2798), .CK(clk), .RN(n4492), .Q(
        \key_mem[8][91] ) );
  DFFRX1 \key_mem_reg[0][59]  ( .D(n1806), .CK(clk), .RN(n4493), .Q(
        \key_mem[0][59] ) );
  DFFRX1 \key_mem_reg[4][59]  ( .D(n2318), .CK(clk), .RN(n4494), .Q(
        \key_mem[4][59] ) );
  DFFRX1 \key_mem_reg[8][59]  ( .D(n2830), .CK(clk), .RN(n4494), .Q(
        \key_mem[8][59] ) );
  DFFRX1 \key_mem_reg[0][27]  ( .D(n1838), .CK(clk), .RN(n4495), .Q(
        \key_mem[0][27] ) );
  DFFRX1 \key_mem_reg[4][27]  ( .D(n2350), .CK(clk), .RN(n4495), .Q(
        \key_mem[4][27] ) );
  DFFRX1 \key_mem_reg[8][27]  ( .D(n2862), .CK(clk), .RN(n4470), .Q(
        \key_mem[8][27] ) );
  DFFRX1 \key_mem_reg[0][126]  ( .D(n1739), .CK(clk), .RN(n4471), .Q(
        \key_mem[0][126] ) );
  DFFRX1 \key_mem_reg[4][126]  ( .D(n2251), .CK(clk), .RN(n4471), .Q(
        \key_mem[4][126] ) );
  DFFRX1 \key_mem_reg[8][126]  ( .D(n2763), .CK(clk), .RN(n4472), .Q(
        \key_mem[8][126] ) );
  DFFRX1 \key_mem_reg[0][94]  ( .D(n1771), .CK(clk), .RN(n4473), .Q(
        \key_mem[0][94] ) );
  DFFRX1 \key_mem_reg[4][94]  ( .D(n2283), .CK(clk), .RN(n4473), .Q(
        \key_mem[4][94] ) );
  DFFRX1 \key_mem_reg[8][94]  ( .D(n2795), .CK(clk), .RN(n4474), .Q(
        \key_mem[8][94] ) );
  DFFRX1 \key_mem_reg[0][62]  ( .D(n1803), .CK(clk), .RN(n4474), .Q(
        \key_mem[0][62] ) );
  DFFRX1 \key_mem_reg[4][62]  ( .D(n2315), .CK(clk), .RN(n4475), .Q(
        \key_mem[4][62] ) );
  DFFRX1 \key_mem_reg[8][62]  ( .D(n2827), .CK(clk), .RN(n4475), .Q(
        \key_mem[8][62] ) );
  DFFRX1 \key_mem_reg[0][30]  ( .D(n1835), .CK(clk), .RN(n4476), .Q(
        \key_mem[0][30] ) );
  DFFRX1 \key_mem_reg[4][30]  ( .D(n2347), .CK(clk), .RN(n4477), .Q(
        \key_mem[4][30] ) );
  DFFRX1 \key_mem_reg[8][30]  ( .D(n2859), .CK(clk), .RN(n4477), .Q(
        \key_mem[8][30] ) );
  DFFRX1 \key_mem_reg[0][125]  ( .D(n1740), .CK(clk), .RN(n4478), .Q(
        \key_mem[0][125] ) );
  DFFRX1 \key_mem_reg[4][125]  ( .D(n2252), .CK(clk), .RN(n4478), .Q(
        \key_mem[4][125] ) );
  DFFRX1 \key_mem_reg[8][125]  ( .D(n2764), .CK(clk), .RN(n4479), .Q(
        \key_mem[8][125] ) );
  DFFRX1 \key_mem_reg[0][93]  ( .D(n1772), .CK(clk), .RN(n4480), .Q(
        \key_mem[0][93] ) );
  DFFRX1 \key_mem_reg[4][93]  ( .D(n2284), .CK(clk), .RN(n4480), .Q(
        \key_mem[4][93] ) );
  DFFRX1 \key_mem_reg[8][93]  ( .D(n2796), .CK(clk), .RN(n4481), .Q(
        \key_mem[8][93] ) );
  DFFRX1 \key_mem_reg[0][61]  ( .D(n1804), .CK(clk), .RN(n4482), .Q(
        \key_mem[0][61] ) );
  DFFRX1 \key_mem_reg[4][61]  ( .D(n2316), .CK(clk), .RN(n4482), .Q(
        \key_mem[4][61] ) );
  DFFRX1 \key_mem_reg[8][61]  ( .D(n2828), .CK(clk), .RN(n4482), .Q(
        \key_mem[8][61] ) );
  DFFRX1 \key_mem_reg[0][29]  ( .D(n1836), .CK(clk), .RN(n4483), .Q(
        \key_mem[0][29] ) );
  DFFRX1 \key_mem_reg[4][29]  ( .D(n2348), .CK(clk), .RN(n4484), .Q(
        \key_mem[4][29] ) );
  DFFRX1 \key_mem_reg[8][29]  ( .D(n2860), .CK(clk), .RN(n4484), .Q(
        \key_mem[8][29] ) );
  DFFRX1 \key_mem_reg[0][124]  ( .D(n1741), .CK(clk), .RN(n4511), .Q(
        \key_mem[0][124] ) );
  DFFRX1 \key_mem_reg[4][124]  ( .D(n2253), .CK(clk), .RN(n4512), .Q(
        \key_mem[4][124] ) );
  DFFRX1 \key_mem_reg[8][124]  ( .D(n2765), .CK(clk), .RN(n4512), .Q(
        \key_mem[8][124] ) );
  DFFRX1 \key_mem_reg[0][92]  ( .D(n1773), .CK(clk), .RN(n4513), .Q(
        \key_mem[0][92] ) );
  DFFRX1 \key_mem_reg[4][92]  ( .D(n2285), .CK(clk), .RN(n4513), .Q(
        \key_mem[4][92] ) );
  DFFRX1 \key_mem_reg[8][92]  ( .D(n2797), .CK(clk), .RN(n4514), .Q(
        \key_mem[8][92] ) );
  DFFRX1 \key_mem_reg[0][60]  ( .D(n1805), .CK(clk), .RN(n4515), .Q(
        \key_mem[0][60] ) );
  DFFRX1 \key_mem_reg[4][60]  ( .D(n2317), .CK(clk), .RN(n4515), .Q(
        \key_mem[4][60] ) );
  DFFRX1 \key_mem_reg[8][60]  ( .D(n2829), .CK(clk), .RN(n4516), .Q(
        \key_mem[8][60] ) );
  DFFRX1 \key_mem_reg[0][28]  ( .D(n1837), .CK(clk), .RN(n4516), .Q(
        \key_mem[0][28] ) );
  DFFRX1 \key_mem_reg[4][28]  ( .D(n2349), .CK(clk), .RN(n4517), .Q(
        \key_mem[4][28] ) );
  DFFRX1 \key_mem_reg[8][28]  ( .D(n2861), .CK(clk), .RN(n4517), .Q(
        \key_mem[8][28] ) );
  DFFRX1 \key_mem_reg[0][121]  ( .D(n1744), .CK(clk), .RN(n4518), .Q(
        \key_mem[0][121] ) );
  DFFRX1 \key_mem_reg[4][121]  ( .D(n2256), .CK(clk), .RN(n4519), .Q(
        \key_mem[4][121] ) );
  DFFRX1 \key_mem_reg[8][121]  ( .D(n2768), .CK(clk), .RN(n4519), .Q(
        \key_mem[8][121] ) );
  DFFRX1 \key_mem_reg[0][89]  ( .D(n1776), .CK(clk), .RN(n4520), .Q(
        \key_mem[0][89] ) );
  DFFRX1 \key_mem_reg[4][89]  ( .D(n2288), .CK(clk), .RN(n4520), .Q(
        \key_mem[4][89] ) );
  DFFRX1 \key_mem_reg[8][89]  ( .D(n2800), .CK(clk), .RN(n4521), .Q(
        \key_mem[8][89] ) );
  DFFRX1 \key_mem_reg[0][57]  ( .D(n1808), .CK(clk), .RN(n4522), .Q(
        \key_mem[0][57] ) );
  DFFRX1 \key_mem_reg[4][57]  ( .D(n2320), .CK(clk), .RN(n4522), .Q(
        \key_mem[4][57] ) );
  DFFRX1 \key_mem_reg[8][57]  ( .D(n2832), .CK(clk), .RN(n4523), .Q(
        \key_mem[8][57] ) );
  DFFRX1 \key_mem_reg[0][25]  ( .D(n1840), .CK(clk), .RN(n4524), .Q(
        \key_mem[0][25] ) );
  DFFRX1 \key_mem_reg[4][25]  ( .D(n2352), .CK(clk), .RN(n4524), .Q(
        \key_mem[4][25] ) );
  DFFRX1 \key_mem_reg[8][25]  ( .D(n2864), .CK(clk), .RN(n4524), .Q(
        \key_mem[8][25] ) );
  DFFRX1 \key_mem_reg[2][119]  ( .D(n2002), .CK(clk), .RN(n4430), .Q(
        \key_mem[2][119] ) );
  DFFRX1 \key_mem_reg[6][119]  ( .D(n2514), .CK(clk), .RN(n4430), .Q(
        \key_mem[6][119] ) );
  DFFRX1 \key_mem_reg[10][119]  ( .D(n3026), .CK(clk), .RN(n4431), .Q(
        \key_mem[10][119] ) );
  DFFRX1 \key_mem_reg[2][118]  ( .D(n2003), .CK(clk), .RN(n4432), .Q(
        \key_mem[2][118] ) );
  DFFRX1 \key_mem_reg[6][118]  ( .D(n2515), .CK(clk), .RN(n4432), .Q(
        \key_mem[6][118] ) );
  DFFRX1 \key_mem_reg[10][118]  ( .D(n3027), .CK(clk), .RN(n4370), .Q(
        \key_mem[10][118] ) );
  DFFRX1 \key_mem_reg[2][117]  ( .D(n2004), .CK(clk), .RN(n4409), .Q(
        \key_mem[2][117] ) );
  DFFRX1 \key_mem_reg[6][117]  ( .D(n2516), .CK(clk), .RN(n4433), .Q(
        \key_mem[6][117] ) );
  DFFRX1 \key_mem_reg[10][117]  ( .D(n3028), .CK(clk), .RN(n4433), .Q(
        \key_mem[10][117] ) );
  DFFRX1 \key_mem_reg[2][116]  ( .D(n2005), .CK(clk), .RN(n4495), .Q(
        \key_mem[2][116] ) );
  DFFRX1 \key_mem_reg[6][116]  ( .D(n2517), .CK(clk), .RN(n4401), .Q(
        \key_mem[6][116] ) );
  DFFRX1 \key_mem_reg[10][116]  ( .D(n3029), .CK(clk), .RN(n4400), .Q(
        \key_mem[10][116] ) );
  DFFRX1 \key_mem_reg[2][115]  ( .D(n2006), .CK(clk), .RN(n4393), .Q(
        \key_mem[2][115] ) );
  DFFRX1 \key_mem_reg[6][115]  ( .D(n2518), .CK(clk), .RN(n4392), .Q(
        \key_mem[6][115] ) );
  DFFRX1 \key_mem_reg[10][115]  ( .D(n3030), .CK(clk), .RN(n4434), .Q(
        \key_mem[10][115] ) );
  DFFRX1 \key_mem_reg[2][114]  ( .D(n2007), .CK(clk), .RN(n4435), .Q(
        \key_mem[2][114] ) );
  DFFRX1 \key_mem_reg[6][114]  ( .D(n2519), .CK(clk), .RN(n4435), .Q(
        \key_mem[6][114] ) );
  DFFRX1 \key_mem_reg[10][114]  ( .D(n3031), .CK(clk), .RN(n4436), .Q(
        \key_mem[10][114] ) );
  DFFRX1 \key_mem_reg[2][113]  ( .D(n2008), .CK(clk), .RN(n4436), .Q(
        \key_mem[2][113] ) );
  DFFRX1 \key_mem_reg[6][113]  ( .D(n2520), .CK(clk), .RN(n4437), .Q(
        \key_mem[6][113] ) );
  DFFRX1 \key_mem_reg[10][113]  ( .D(n3032), .CK(clk), .RN(n4437), .Q(
        \key_mem[10][113] ) );
  DFFRX1 \key_mem_reg[2][112]  ( .D(n2009), .CK(clk), .RN(n4438), .Q(
        \key_mem[2][112] ) );
  DFFRX1 \key_mem_reg[6][112]  ( .D(n2521), .CK(clk), .RN(n4439), .Q(
        \key_mem[6][112] ) );
  DFFRX1 \key_mem_reg[10][112]  ( .D(n3033), .CK(clk), .RN(n4439), .Q(
        \key_mem[10][112] ) );
  DFFRX1 \key_mem_reg[2][111]  ( .D(n2010), .CK(clk), .RN(n4440), .Q(
        \key_mem[2][111] ) );
  DFFRX1 \key_mem_reg[6][111]  ( .D(n2522), .CK(clk), .RN(n4417), .Q(
        \key_mem[6][111] ) );
  DFFRX1 \key_mem_reg[10][111]  ( .D(n3034), .CK(clk), .RN(n4418), .Q(
        \key_mem[10][111] ) );
  DFFRX1 \key_mem_reg[2][110]  ( .D(n2011), .CK(clk), .RN(n4418), .Q(
        \key_mem[2][110] ) );
  DFFRX1 \key_mem_reg[6][110]  ( .D(n2523), .CK(clk), .RN(n4436), .Q(
        \key_mem[6][110] ) );
  DFFRX1 \key_mem_reg[10][110]  ( .D(n3035), .CK(clk), .RN(n4434), .Q(
        \key_mem[10][110] ) );
  DFFRX1 \key_mem_reg[2][109]  ( .D(n2012), .CK(clk), .RN(n4419), .Q(
        \key_mem[2][109] ) );
  DFFRX1 \key_mem_reg[6][109]  ( .D(n2524), .CK(clk), .RN(n4420), .Q(
        \key_mem[6][109] ) );
  DFFRX1 \key_mem_reg[10][109]  ( .D(n3036), .CK(clk), .RN(n4420), .Q(
        \key_mem[10][109] ) );
  DFFRX1 \key_mem_reg[2][108]  ( .D(n2013), .CK(clk), .RN(n4421), .Q(
        \key_mem[2][108] ) );
  DFFRX1 \key_mem_reg[6][108]  ( .D(n2525), .CK(clk), .RN(n4421), .Q(
        \key_mem[6][108] ) );
  DFFRX1 \key_mem_reg[10][108]  ( .D(n3037), .CK(clk), .RN(n4422), .Q(
        \key_mem[10][108] ) );
  DFFRX1 \key_mem_reg[2][106]  ( .D(n2015), .CK(clk), .RN(n4423), .Q(
        \key_mem[2][106] ) );
  DFFRX1 \key_mem_reg[6][106]  ( .D(n2527), .CK(clk), .RN(n4423), .Q(
        \key_mem[6][106] ) );
  DFFRX1 \key_mem_reg[10][106]  ( .D(n3039), .CK(clk), .RN(n4424), .Q(
        \key_mem[10][106] ) );
  DFFRX1 \key_mem_reg[2][105]  ( .D(n2016), .CK(clk), .RN(n4424), .Q(
        \key_mem[2][105] ) );
  DFFRX1 \key_mem_reg[6][105]  ( .D(n2528), .CK(clk), .RN(n4425), .Q(
        \key_mem[6][105] ) );
  DFFRX1 \key_mem_reg[10][105]  ( .D(n3040), .CK(clk), .RN(n4425), .Q(
        \key_mem[10][105] ) );
  DFFRX1 \key_mem_reg[2][104]  ( .D(n2017), .CK(clk), .RN(n4426), .Q(
        \key_mem[2][104] ) );
  DFFRX1 \key_mem_reg[6][104]  ( .D(n2529), .CK(clk), .RN(n4427), .Q(
        \key_mem[6][104] ) );
  DFFRX1 \key_mem_reg[10][104]  ( .D(n3041), .CK(clk), .RN(n4427), .Q(
        \key_mem[10][104] ) );
  DFFRX1 \key_mem_reg[2][103]  ( .D(n2018), .CK(clk), .RN(n4428), .Q(
        \key_mem[2][103] ) );
  DFFRX1 \key_mem_reg[6][103]  ( .D(n2530), .CK(clk), .RN(n4428), .Q(
        \key_mem[6][103] ) );
  DFFRX1 \key_mem_reg[10][103]  ( .D(n3042), .CK(clk), .RN(n4429), .Q(
        \key_mem[10][103] ) );
  DFFRX1 \key_mem_reg[2][102]  ( .D(n2019), .CK(clk), .RN(n4456), .Q(
        \key_mem[2][102] ) );
  DFFRX1 \key_mem_reg[6][102]  ( .D(n2531), .CK(clk), .RN(n4456), .Q(
        \key_mem[6][102] ) );
  DFFRX1 \key_mem_reg[10][102]  ( .D(n3043), .CK(clk), .RN(n4457), .Q(
        \key_mem[10][102] ) );
  DFFRX1 \key_mem_reg[2][101]  ( .D(n2020), .CK(clk), .RN(n4457), .Q(
        \key_mem[2][101] ) );
  DFFRX1 \key_mem_reg[6][101]  ( .D(n2532), .CK(clk), .RN(n4458), .Q(
        \key_mem[6][101] ) );
  DFFRX1 \key_mem_reg[10][101]  ( .D(n3044), .CK(clk), .RN(n4458), .Q(
        \key_mem[10][101] ) );
  DFFRX1 \key_mem_reg[2][100]  ( .D(n2021), .CK(clk), .RN(n4459), .Q(
        \key_mem[2][100] ) );
  DFFRX1 \key_mem_reg[6][100]  ( .D(n2533), .CK(clk), .RN(n4460), .Q(
        \key_mem[6][100] ) );
  DFFRX1 \key_mem_reg[10][100]  ( .D(n3045), .CK(clk), .RN(n4460), .Q(
        \key_mem[10][100] ) );
  DFFRX1 \key_mem_reg[2][99]  ( .D(n2022), .CK(clk), .RN(n4471), .Q(
        \key_mem[2][99] ) );
  DFFRX1 \key_mem_reg[6][99]  ( .D(n2534), .CK(clk), .RN(n4470), .Q(
        \key_mem[6][99] ) );
  DFFRX1 \key_mem_reg[10][99]  ( .D(n3046), .CK(clk), .RN(n4461), .Q(
        \key_mem[10][99] ) );
  DFFRX1 \key_mem_reg[2][98]  ( .D(n2023), .CK(clk), .RN(n4462), .Q(
        \key_mem[2][98] ) );
  DFFRX1 \key_mem_reg[6][98]  ( .D(n2535), .CK(clk), .RN(n4462), .Q(
        \key_mem[6][98] ) );
  DFFRX1 \key_mem_reg[10][98]  ( .D(n3047), .CK(clk), .RN(n4463), .Q(
        \key_mem[10][98] ) );
  DFFRX1 \key_mem_reg[2][97]  ( .D(n2024), .CK(clk), .RN(n4464), .Q(
        \key_mem[2][97] ) );
  DFFRX1 \key_mem_reg[6][97]  ( .D(n2536), .CK(clk), .RN(n4464), .Q(
        \key_mem[6][97] ) );
  DFFRX1 \key_mem_reg[10][97]  ( .D(n3048), .CK(clk), .RN(n4465), .Q(
        \key_mem[10][97] ) );
  DFFRX1 \key_mem_reg[2][96]  ( .D(n2025), .CK(clk), .RN(n4465), .Q(
        \key_mem[2][96] ) );
  DFFRX1 \key_mem_reg[6][96]  ( .D(n2537), .CK(clk), .RN(n4466), .Q(
        \key_mem[6][96] ) );
  DFFRX1 \key_mem_reg[10][96]  ( .D(n3049), .CK(clk), .RN(n4466), .Q(
        \key_mem[10][96] ) );
  DFFRX1 \key_mem_reg[2][87]  ( .D(n2034), .CK(clk), .RN(n4467), .Q(
        \key_mem[2][87] ) );
  DFFRX1 \key_mem_reg[6][87]  ( .D(n2546), .CK(clk), .RN(n4468), .Q(
        \key_mem[6][87] ) );
  DFFRX1 \key_mem_reg[10][87]  ( .D(n3058), .CK(clk), .RN(n4468), .Q(
        \key_mem[10][87] ) );
  DFFRX1 \key_mem_reg[2][86]  ( .D(n2035), .CK(clk), .RN(n4469), .Q(
        \key_mem[2][86] ) );
  DFFRX1 \key_mem_reg[6][86]  ( .D(n2547), .CK(clk), .RN(n4469), .Q(
        \key_mem[6][86] ) );
  DFFRX1 \key_mem_reg[10][86]  ( .D(n3059), .CK(clk), .RN(n4441), .Q(
        \key_mem[10][86] ) );
  DFFRX1 \key_mem_reg[2][85]  ( .D(n2036), .CK(clk), .RN(n4441), .Q(
        \key_mem[2][85] ) );
  DFFRX1 \key_mem_reg[6][85]  ( .D(n2548), .CK(clk), .RN(n4442), .Q(
        \key_mem[6][85] ) );
  DFFRX1 \key_mem_reg[10][85]  ( .D(n3060), .CK(clk), .RN(n4442), .Q(
        \key_mem[10][85] ) );
  DFFRX1 \key_mem_reg[2][84]  ( .D(n2037), .CK(clk), .RN(n4443), .Q(
        \key_mem[2][84] ) );
  DFFRX1 \key_mem_reg[6][84]  ( .D(n2549), .CK(clk), .RN(n4444), .Q(
        \key_mem[6][84] ) );
  DFFRX1 \key_mem_reg[10][84]  ( .D(n3061), .CK(clk), .RN(n4444), .Q(
        \key_mem[10][84] ) );
  DFFRX1 \key_mem_reg[2][83]  ( .D(n2038), .CK(clk), .RN(n4445), .Q(
        \key_mem[2][83] ) );
  DFFRX1 \key_mem_reg[6][83]  ( .D(n2550), .CK(clk), .RN(n4445), .Q(
        \key_mem[6][83] ) );
  DFFRX1 \key_mem_reg[10][83]  ( .D(n3062), .CK(clk), .RN(n4446), .Q(
        \key_mem[10][83] ) );
  DFFRX1 \key_mem_reg[2][82]  ( .D(n2039), .CK(clk), .RN(n4447), .Q(
        \key_mem[2][82] ) );
  DFFRX1 \key_mem_reg[6][82]  ( .D(n2551), .CK(clk), .RN(n4447), .Q(
        \key_mem[6][82] ) );
  DFFRX1 \key_mem_reg[10][82]  ( .D(n3063), .CK(clk), .RN(n4448), .Q(
        \key_mem[10][82] ) );
  DFFRX1 \key_mem_reg[2][81]  ( .D(n2040), .CK(clk), .RN(n4448), .Q(
        \key_mem[2][81] ) );
  DFFRX1 \key_mem_reg[6][81]  ( .D(n2552), .CK(clk), .RN(n4449), .Q(
        \key_mem[6][81] ) );
  DFFRX1 \key_mem_reg[10][81]  ( .D(n3064), .CK(clk), .RN(n4449), .Q(
        \key_mem[10][81] ) );
  DFFRX1 \key_mem_reg[2][80]  ( .D(n2041), .CK(clk), .RN(n4450), .Q(
        \key_mem[2][80] ) );
  DFFRX1 \key_mem_reg[6][80]  ( .D(n2553), .CK(clk), .RN(n4451), .Q(
        \key_mem[6][80] ) );
  DFFRX1 \key_mem_reg[10][80]  ( .D(n3065), .CK(clk), .RN(n4451), .Q(
        \key_mem[10][80] ) );
  DFFRX1 \key_mem_reg[2][79]  ( .D(n2042), .CK(clk), .RN(n4452), .Q(
        \key_mem[2][79] ) );
  DFFRX1 \key_mem_reg[6][79]  ( .D(n2554), .CK(clk), .RN(n4452), .Q(
        \key_mem[6][79] ) );
  DFFRX1 \key_mem_reg[10][79]  ( .D(n3066), .CK(clk), .RN(n4453), .Q(
        \key_mem[10][79] ) );
  DFFRX1 \key_mem_reg[2][78]  ( .D(n2043), .CK(clk), .RN(n4454), .Q(
        \key_mem[2][78] ) );
  DFFRX1 \key_mem_reg[6][78]  ( .D(n2555), .CK(clk), .RN(n4454), .Q(
        \key_mem[6][78] ) );
  DFFRX1 \key_mem_reg[10][78]  ( .D(n3067), .CK(clk), .RN(n4455), .Q(
        \key_mem[10][78] ) );
  DFFRX1 \key_mem_reg[2][77]  ( .D(n2044), .CK(clk), .RN(n4455), .Q(
        \key_mem[2][77] ) );
  DFFRX1 \key_mem_reg[6][77]  ( .D(n2556), .CK(clk), .RN(n4373), .Q(
        \key_mem[6][77] ) );
  DFFRX1 \key_mem_reg[10][77]  ( .D(n3068), .CK(clk), .RN(n4373), .Q(
        \key_mem[10][77] ) );
  DFFRX1 \key_mem_reg[2][76]  ( .D(n2045), .CK(clk), .RN(n4374), .Q(
        \key_mem[2][76] ) );
  DFFRX1 \key_mem_reg[6][76]  ( .D(n2557), .CK(clk), .RN(n4375), .Q(
        \key_mem[6][76] ) );
  DFFRX1 \key_mem_reg[10][76]  ( .D(n3069), .CK(clk), .RN(n4375), .Q(
        \key_mem[10][76] ) );
  DFFRX1 \key_mem_reg[2][75]  ( .D(n2046), .CK(clk), .RN(n4376), .Q(
        \key_mem[2][75] ) );
  DFFRX1 \key_mem_reg[6][75]  ( .D(n2558), .CK(clk), .RN(n4376), .Q(
        \key_mem[6][75] ) );
  DFFRX1 \key_mem_reg[10][75]  ( .D(n3070), .CK(clk), .RN(n4377), .Q(
        \key_mem[10][75] ) );
  DFFRX1 \key_mem_reg[2][74]  ( .D(n2047), .CK(clk), .RN(n4378), .Q(
        \key_mem[2][74] ) );
  DFFRX1 \key_mem_reg[6][74]  ( .D(n2559), .CK(clk), .RN(n4378), .Q(
        \key_mem[6][74] ) );
  DFFRX1 \key_mem_reg[10][74]  ( .D(n3071), .CK(clk), .RN(n4379), .Q(
        \key_mem[10][74] ) );
  DFFRX1 \key_mem_reg[2][73]  ( .D(n2048), .CK(clk), .RN(n4379), .Q(
        \key_mem[2][73] ) );
  DFFRX1 \key_mem_reg[6][73]  ( .D(n2560), .CK(clk), .RN(n4380), .Q(
        \key_mem[6][73] ) );
  DFFRX1 \key_mem_reg[10][73]  ( .D(n3072), .CK(clk), .RN(n4381), .Q(
        \key_mem[10][73] ) );
  DFFRX1 \key_mem_reg[2][72]  ( .D(n2049), .CK(clk), .RN(n4381), .Q(
        \key_mem[2][72] ) );
  DFFRX1 \key_mem_reg[6][72]  ( .D(n2561), .CK(clk), .RN(n4382), .Q(
        \key_mem[6][72] ) );
  DFFRX1 \key_mem_reg[10][72]  ( .D(n3073), .CK(clk), .RN(n4382), .Q(
        \key_mem[10][72] ) );
  DFFRX1 \key_mem_reg[2][71]  ( .D(n2050), .CK(clk), .RN(n4383), .Q(
        \key_mem[2][71] ) );
  DFFRX1 \key_mem_reg[6][71]  ( .D(n2562), .CK(clk), .RN(n4384), .Q(
        \key_mem[6][71] ) );
  DFFRX1 \key_mem_reg[10][71]  ( .D(n3074), .CK(clk), .RN(n4384), .Q(
        \key_mem[10][71] ) );
  DFFRX1 \key_mem_reg[2][70]  ( .D(n2051), .CK(clk), .RN(n4385), .Q(
        \key_mem[2][70] ) );
  DFFRX1 \key_mem_reg[6][70]  ( .D(n2563), .CK(clk), .RN(n4385), .Q(
        \key_mem[6][70] ) );
  DFFRX1 \key_mem_reg[10][70]  ( .D(n3075), .CK(clk), .RN(n4386), .Q(
        \key_mem[10][70] ) );
  DFFRX1 \key_mem_reg[2][69]  ( .D(n2052), .CK(clk), .RN(n4387), .Q(
        \key_mem[2][69] ) );
  DFFRX1 \key_mem_reg[6][69]  ( .D(n2564), .CK(clk), .RN(n4387), .Q(
        \key_mem[6][69] ) );
  DFFRX1 \key_mem_reg[10][69]  ( .D(n3076), .CK(clk), .RN(n4388), .Q(
        \key_mem[10][69] ) );
  DFFRX1 \key_mem_reg[2][68]  ( .D(n2053), .CK(clk), .RN(n4502), .Q(
        \key_mem[2][68] ) );
  DFFRX1 \key_mem_reg[6][68]  ( .D(n2565), .CK(clk), .RN(n4392), .Q(
        \key_mem[6][68] ) );
  DFFRX1 \key_mem_reg[10][68]  ( .D(n3077), .CK(clk), .RN(n4423), .Q(
        \key_mem[10][68] ) );
  DFFRX1 \key_mem_reg[2][67]  ( .D(n2054), .CK(clk), .RN(n4386), .Q(
        \key_mem[2][67] ) );
  DFFRX1 \key_mem_reg[6][67]  ( .D(n2566), .CK(clk), .RN(n4385), .Q(
        \key_mem[6][67] ) );
  DFFRX1 \key_mem_reg[10][67]  ( .D(n3078), .CK(clk), .RN(n4373), .Q(
        \key_mem[10][67] ) );
  DFFRX1 \key_mem_reg[2][66]  ( .D(n2055), .CK(clk), .RN(n4403), .Q(
        \key_mem[2][66] ) );
  DFFRX1 \key_mem_reg[6][66]  ( .D(n2567), .CK(clk), .RN(n4402), .Q(
        \key_mem[6][66] ) );
  DFFRX1 \key_mem_reg[10][66]  ( .D(n3079), .CK(clk), .RN(n4395), .Q(
        \key_mem[10][66] ) );
  DFFRX1 \key_mem_reg[2][65]  ( .D(n2056), .CK(clk), .RN(n4396), .Q(
        \key_mem[2][65] ) );
  DFFRX1 \key_mem_reg[6][65]  ( .D(n2568), .CK(clk), .RN(n4451), .Q(
        \key_mem[6][65] ) );
  DFFRX1 \key_mem_reg[10][65]  ( .D(n3080), .CK(clk), .RN(n4452), .Q(
        \key_mem[10][65] ) );
  DFFRX1 \key_mem_reg[2][64]  ( .D(n2057), .CK(clk), .RN(n4446), .Q(
        \key_mem[2][64] ) );
  DFFRX1 \key_mem_reg[6][64]  ( .D(n2569), .CK(clk), .RN(n4450), .Q(
        \key_mem[6][64] ) );
  DFFRX1 \key_mem_reg[10][64]  ( .D(n3081), .CK(clk), .RN(n4460), .Q(
        \key_mem[10][64] ) );
  DFFRX1 \key_mem_reg[2][55]  ( .D(n2066), .CK(clk), .RN(n4538), .Q(
        \key_mem[2][55] ) );
  DFFRX1 \key_mem_reg[6][55]  ( .D(n2578), .CK(clk), .RN(n4552), .Q(
        \key_mem[6][55] ) );
  DFFRX1 \key_mem_reg[10][55]  ( .D(n3090), .CK(clk), .RN(n4551), .Q(
        \key_mem[10][55] ) );
  DFFRX1 \key_mem_reg[2][54]  ( .D(n2067), .CK(clk), .RN(n4538), .Q(
        \key_mem[2][54] ) );
  DFFRX1 \key_mem_reg[6][54]  ( .D(n2579), .CK(clk), .RN(n4537), .Q(
        \key_mem[6][54] ) );
  DFFRX1 \key_mem_reg[10][54]  ( .D(n3091), .CK(clk), .RN(n4370), .Q(
        \key_mem[10][54] ) );
  DFFRX1 \key_mem_reg[2][53]  ( .D(n2068), .CK(clk), .RN(n4371), .Q(
        \key_mem[2][53] ) );
  DFFRX1 \key_mem_reg[6][53]  ( .D(n2580), .CK(clk), .RN(n4371), .Q(
        \key_mem[6][53] ) );
  DFFRX1 \key_mem_reg[10][53]  ( .D(n3092), .CK(clk), .RN(n4372), .Q(
        \key_mem[10][53] ) );
  DFFRX1 \key_mem_reg[2][52]  ( .D(n2069), .CK(clk), .RN(n4372), .Q(
        \key_mem[2][52] ) );
  DFFRX1 \key_mem_reg[6][52]  ( .D(n2581), .CK(clk), .RN(n4410), .Q(
        \key_mem[6][52] ) );
  DFFRX1 \key_mem_reg[10][52]  ( .D(n3093), .CK(clk), .RN(n4403), .Q(
        \key_mem[10][52] ) );
  DFFRX1 \key_mem_reg[2][51]  ( .D(n2070), .CK(clk), .RN(n4404), .Q(
        \key_mem[2][51] ) );
  DFFRX1 \key_mem_reg[6][51]  ( .D(n2582), .CK(clk), .RN(n4405), .Q(
        \key_mem[6][51] ) );
  DFFRX1 \key_mem_reg[10][51]  ( .D(n3094), .CK(clk), .RN(n4405), .Q(
        \key_mem[10][51] ) );
  DFFRX1 \key_mem_reg[2][50]  ( .D(n2071), .CK(clk), .RN(n4406), .Q(
        \key_mem[2][50] ) );
  DFFRX1 \key_mem_reg[6][50]  ( .D(n2583), .CK(clk), .RN(n4406), .Q(
        \key_mem[6][50] ) );
  DFFRX1 \key_mem_reg[10][50]  ( .D(n3095), .CK(clk), .RN(n4407), .Q(
        \key_mem[10][50] ) );
  DFFRX1 \key_mem_reg[2][49]  ( .D(n2072), .CK(clk), .RN(n4408), .Q(
        \key_mem[2][49] ) );
  DFFRX1 \key_mem_reg[6][49]  ( .D(n2584), .CK(clk), .RN(n4408), .Q(
        \key_mem[6][49] ) );
  DFFRX1 \key_mem_reg[10][49]  ( .D(n3096), .CK(clk), .RN(n4409), .Q(
        \key_mem[10][49] ) );
  DFFRX1 \key_mem_reg[2][47]  ( .D(n2074), .CK(clk), .RN(n4411), .Q(
        \key_mem[2][47] ) );
  DFFRX1 \key_mem_reg[6][47]  ( .D(n2586), .CK(clk), .RN(n4412), .Q(
        \key_mem[6][47] ) );
  DFFRX1 \key_mem_reg[10][47]  ( .D(n3098), .CK(clk), .RN(n4412), .Q(
        \key_mem[10][47] ) );
  DFFRX1 \key_mem_reg[2][46]  ( .D(n2075), .CK(clk), .RN(n4413), .Q(
        \key_mem[2][46] ) );
  DFFRX1 \key_mem_reg[6][46]  ( .D(n2587), .CK(clk), .RN(n4377), .Q(
        \key_mem[6][46] ) );
  DFFRX1 \key_mem_reg[10][46]  ( .D(n3099), .CK(clk), .RN(n4387), .Q(
        \key_mem[10][46] ) );
  DFFRX1 \key_mem_reg[2][45]  ( .D(n2076), .CK(clk), .RN(n4414), .Q(
        \key_mem[2][45] ) );
  DFFRX1 \key_mem_reg[6][45]  ( .D(n2588), .CK(clk), .RN(n4414), .Q(
        \key_mem[6][45] ) );
  DFFRX1 \key_mem_reg[10][45]  ( .D(n3100), .CK(clk), .RN(n4415), .Q(
        \key_mem[10][45] ) );
  DFFRX1 \key_mem_reg[2][44]  ( .D(n2077), .CK(clk), .RN(n4416), .Q(
        \key_mem[2][44] ) );
  DFFRX1 \key_mem_reg[6][44]  ( .D(n2589), .CK(clk), .RN(n4416), .Q(
        \key_mem[6][44] ) );
  DFFRX1 \key_mem_reg[10][44]  ( .D(n3101), .CK(clk), .RN(n4417), .Q(
        \key_mem[10][44] ) );
  DFFRX1 \key_mem_reg[2][43]  ( .D(n2078), .CK(clk), .RN(n4388), .Q(
        \key_mem[2][43] ) );
  DFFRX1 \key_mem_reg[6][43]  ( .D(n2590), .CK(clk), .RN(n4389), .Q(
        \key_mem[6][43] ) );
  DFFRX1 \key_mem_reg[10][43]  ( .D(n3102), .CK(clk), .RN(n4389), .Q(
        \key_mem[10][43] ) );
  DFFRX1 \key_mem_reg[2][42]  ( .D(n2079), .CK(clk), .RN(n4390), .Q(
        \key_mem[2][42] ) );
  DFFRX1 \key_mem_reg[6][42]  ( .D(n2591), .CK(clk), .RN(n4390), .Q(
        \key_mem[6][42] ) );
  DFFRX1 \key_mem_reg[10][42]  ( .D(n3103), .CK(clk), .RN(n4391), .Q(
        \key_mem[10][42] ) );
  DFFRX1 \key_mem_reg[2][41]  ( .D(n2080), .CK(clk), .RN(n4392), .Q(
        \key_mem[2][41] ) );
  DFFRX1 \key_mem_reg[6][41]  ( .D(n2592), .CK(clk), .RN(n4392), .Q(
        \key_mem[6][41] ) );
  DFFRX1 \key_mem_reg[10][41]  ( .D(n3104), .CK(clk), .RN(n4393), .Q(
        \key_mem[10][41] ) );
  DFFRX1 \key_mem_reg[2][40]  ( .D(n2081), .CK(clk), .RN(n4393), .Q(
        \key_mem[2][40] ) );
  DFFRX1 \key_mem_reg[6][40]  ( .D(n2593), .CK(clk), .RN(n4394), .Q(
        \key_mem[6][40] ) );
  DFFRX1 \key_mem_reg[10][40]  ( .D(n3105), .CK(clk), .RN(n4394), .Q(
        \key_mem[10][40] ) );
  DFFRX1 \key_mem_reg[2][39]  ( .D(n2082), .CK(clk), .RN(n4395), .Q(
        \key_mem[2][39] ) );
  DFFRX1 \key_mem_reg[6][39]  ( .D(n2594), .CK(clk), .RN(n4396), .Q(
        \key_mem[6][39] ) );
  DFFRX1 \key_mem_reg[10][39]  ( .D(n3106), .CK(clk), .RN(n4396), .Q(
        \key_mem[10][39] ) );
  DFFRX1 \key_mem_reg[2][38]  ( .D(n2083), .CK(clk), .RN(n4397), .Q(
        \key_mem[2][38] ) );
  DFFRX1 \key_mem_reg[6][38]  ( .D(n2595), .CK(clk), .RN(n4397), .Q(
        \key_mem[6][38] ) );
  DFFRX1 \key_mem_reg[10][38]  ( .D(n3107), .CK(clk), .RN(n4398), .Q(
        \key_mem[10][38] ) );
  DFFRX1 \key_mem_reg[2][37]  ( .D(n2084), .CK(clk), .RN(n4399), .Q(
        \key_mem[2][37] ) );
  DFFRX1 \key_mem_reg[6][37]  ( .D(n2596), .CK(clk), .RN(n4399), .Q(
        \key_mem[6][37] ) );
  DFFRX1 \key_mem_reg[10][37]  ( .D(n3108), .CK(clk), .RN(n4400), .Q(
        \key_mem[10][37] ) );
  DFFRX1 \key_mem_reg[2][36]  ( .D(n2085), .CK(clk), .RN(n4400), .Q(
        \key_mem[2][36] ) );
  DFFRX1 \key_mem_reg[6][36]  ( .D(n2597), .CK(clk), .RN(n4401), .Q(
        \key_mem[6][36] ) );
  DFFRX1 \key_mem_reg[10][36]  ( .D(n3109), .CK(clk), .RN(n4401), .Q(
        \key_mem[10][36] ) );
  DFFRX1 \key_mem_reg[2][35]  ( .D(n2086), .CK(clk), .RN(n4402), .Q(
        \key_mem[2][35] ) );
  DFFRX1 \key_mem_reg[6][35]  ( .D(n2598), .CK(clk), .RN(n4403), .Q(
        \key_mem[6][35] ) );
  DFFRX1 \key_mem_reg[10][35]  ( .D(n3110), .CK(clk), .RN(n4554), .Q(
        \key_mem[10][35] ) );
  DFFRX1 \key_mem_reg[2][34]  ( .D(n2087), .CK(clk), .RN(n4542), .Q(
        \key_mem[2][34] ) );
  DFFRX1 \key_mem_reg[6][34]  ( .D(n2599), .CK(clk), .RN(n4542), .Q(
        \key_mem[6][34] ) );
  DFFRX1 \key_mem_reg[10][34]  ( .D(n3111), .CK(clk), .RN(n4543), .Q(
        \key_mem[10][34] ) );
  DFFRX1 \key_mem_reg[2][33]  ( .D(n2088), .CK(clk), .RN(n4544), .Q(
        \key_mem[2][33] ) );
  DFFRX1 \key_mem_reg[6][33]  ( .D(n2600), .CK(clk), .RN(n4544), .Q(
        \key_mem[6][33] ) );
  DFFRX1 \key_mem_reg[10][33]  ( .D(n3112), .CK(clk), .RN(n4545), .Q(
        \key_mem[10][33] ) );
  DFFRX1 \key_mem_reg[2][32]  ( .D(n2089), .CK(clk), .RN(n4545), .Q(
        \key_mem[2][32] ) );
  DFFRX1 \key_mem_reg[6][32]  ( .D(n2601), .CK(clk), .RN(n4546), .Q(
        \key_mem[6][32] ) );
  DFFRX1 \key_mem_reg[10][32]  ( .D(n3113), .CK(clk), .RN(n4546), .Q(
        \key_mem[10][32] ) );
  DFFRX1 \key_mem_reg[2][23]  ( .D(n2098), .CK(clk), .RN(n4547), .Q(
        \key_mem[2][23] ) );
  DFFRX1 \key_mem_reg[6][23]  ( .D(n2610), .CK(clk), .RN(n4548), .Q(
        \key_mem[6][23] ) );
  DFFRX1 \key_mem_reg[10][23]  ( .D(n3122), .CK(clk), .RN(n4548), .Q(
        \key_mem[10][23] ) );
  DFFRX1 \key_mem_reg[2][22]  ( .D(n2099), .CK(clk), .RN(n4549), .Q(
        \key_mem[2][22] ) );
  DFFRX1 \key_mem_reg[6][22]  ( .D(n2611), .CK(clk), .RN(n4549), .Q(
        \key_mem[6][22] ) );
  DFFRX1 \key_mem_reg[10][22]  ( .D(n3123), .CK(clk), .RN(n4550), .Q(
        \key_mem[10][22] ) );
  DFFRX1 \key_mem_reg[2][21]  ( .D(n2100), .CK(clk), .RN(n4551), .Q(
        \key_mem[2][21] ) );
  DFFRX1 \key_mem_reg[6][21]  ( .D(n2612), .CK(clk), .RN(n4551), .Q(
        \key_mem[6][21] ) );
  DFFRX1 \key_mem_reg[10][21]  ( .D(n3124), .CK(clk), .RN(n4552), .Q(
        \key_mem[10][21] ) );
  DFFRX1 \key_mem_reg[2][20]  ( .D(n2101), .CK(clk), .RN(n4552), .Q(
        \key_mem[2][20] ) );
  DFFRX1 \key_mem_reg[6][20]  ( .D(n2613), .CK(clk), .RN(n4553), .Q(
        \key_mem[6][20] ) );
  DFFRX1 \key_mem_reg[10][20]  ( .D(n3125), .CK(clk), .RN(n4553), .Q(
        \key_mem[10][20] ) );
  DFFRX1 \key_mem_reg[2][18]  ( .D(n2103), .CK(clk), .RN(n4554), .Q(
        \key_mem[2][18] ) );
  DFFRX1 \key_mem_reg[6][18]  ( .D(n2615), .CK(clk), .RN(n4526), .Q(
        \key_mem[6][18] ) );
  DFFRX1 \key_mem_reg[10][18]  ( .D(n3127), .CK(clk), .RN(n4527), .Q(
        \key_mem[10][18] ) );
  DFFRX1 \key_mem_reg[2][17]  ( .D(n2104), .CK(clk), .RN(n4527), .Q(
        \key_mem[2][17] ) );
  DFFRX1 \key_mem_reg[6][17]  ( .D(n2616), .CK(clk), .RN(n4528), .Q(
        \key_mem[6][17] ) );
  DFFRX1 \key_mem_reg[10][17]  ( .D(n3128), .CK(clk), .RN(n4528), .Q(
        \key_mem[10][17] ) );
  DFFRX1 \key_mem_reg[2][16]  ( .D(n2105), .CK(clk), .RN(n4529), .Q(
        \key_mem[2][16] ) );
  DFFRX1 \key_mem_reg[6][16]  ( .D(n2617), .CK(clk), .RN(n4530), .Q(
        \key_mem[6][16] ) );
  DFFRX1 \key_mem_reg[10][16]  ( .D(n3129), .CK(clk), .RN(n4530), .Q(
        \key_mem[10][16] ) );
  DFFRX1 \key_mem_reg[2][15]  ( .D(n2106), .CK(clk), .RN(n4531), .Q(
        \key_mem[2][15] ) );
  DFFRX1 \key_mem_reg[6][15]  ( .D(n2618), .CK(clk), .RN(n4531), .Q(
        \key_mem[6][15] ) );
  DFFRX1 \key_mem_reg[10][15]  ( .D(n3130), .CK(clk), .RN(n4532), .Q(
        \key_mem[10][15] ) );
  DFFRX1 \key_mem_reg[2][14]  ( .D(n2107), .CK(clk), .RN(n4533), .Q(
        \key_mem[2][14] ) );
  DFFRX1 \key_mem_reg[6][14]  ( .D(n2619), .CK(clk), .RN(n4533), .Q(
        \key_mem[6][14] ) );
  DFFRX1 \key_mem_reg[10][14]  ( .D(n3131), .CK(clk), .RN(n4534), .Q(
        \key_mem[10][14] ) );
  DFFRX1 \key_mem_reg[2][13]  ( .D(n2108), .CK(clk), .RN(n4535), .Q(
        \key_mem[2][13] ) );
  DFFRX1 \key_mem_reg[6][13]  ( .D(n2620), .CK(clk), .RN(n4535), .Q(
        \key_mem[6][13] ) );
  DFFRX1 \key_mem_reg[10][13]  ( .D(n3132), .CK(clk), .RN(n4536), .Q(
        \key_mem[10][13] ) );
  DFFRX1 \key_mem_reg[2][12]  ( .D(n2109), .CK(clk), .RN(n4536), .Q(
        \key_mem[2][12] ) );
  DFFRX1 \key_mem_reg[6][12]  ( .D(n2621), .CK(clk), .RN(n4537), .Q(
        \key_mem[6][12] ) );
  DFFRX1 \key_mem_reg[10][12]  ( .D(n3133), .CK(clk), .RN(n4537), .Q(
        \key_mem[10][12] ) );
  DFFRX1 \key_mem_reg[2][11]  ( .D(n2110), .CK(clk), .RN(n4538), .Q(
        \key_mem[2][11] ) );
  DFFRX1 \key_mem_reg[6][11]  ( .D(n2622), .CK(clk), .RN(n4539), .Q(
        \key_mem[6][11] ) );
  DFFRX1 \key_mem_reg[10][11]  ( .D(n3134), .CK(clk), .RN(n4539), .Q(
        \key_mem[10][11] ) );
  DFFRX1 \key_mem_reg[2][10]  ( .D(n2111), .CK(clk), .RN(n4540), .Q(
        \key_mem[2][10] ) );
  DFFRX1 \key_mem_reg[6][10]  ( .D(n2623), .CK(clk), .RN(n4540), .Q(
        \key_mem[6][10] ) );
  DFFRX1 \key_mem_reg[10][10]  ( .D(n3135), .CK(clk), .RN(n4541), .Q(
        \key_mem[10][10] ) );
  DFFRX1 \key_mem_reg[2][9]  ( .D(n2112), .CK(clk), .RN(n4533), .Q(
        \key_mem[2][9] ) );
  DFFRX1 \key_mem_reg[6][9]  ( .D(n2624), .CK(clk), .RN(n4532), .Q(
        \key_mem[6][9] ) );
  DFFRX1 \key_mem_reg[10][9]  ( .D(n3136), .CK(clk), .RN(n4528), .Q(
        \key_mem[10][9] ) );
  DFFRX1 \key_mem_reg[2][8]  ( .D(n2113), .CK(clk), .RN(n4523), .Q(
        \key_mem[2][8] ) );
  DFFRX1 \key_mem_reg[6][8]  ( .D(n2625), .CK(clk), .RN(n4495), .Q(
        \key_mem[6][8] ) );
  DFFRX1 \key_mem_reg[10][8]  ( .D(n3137), .CK(clk), .RN(n4520), .Q(
        \key_mem[10][8] ) );
  DFFRX1 \key_mem_reg[2][7]  ( .D(n2114), .CK(clk), .RN(n4559), .Q(
        \key_mem[2][7] ) );
  DFFRX1 \key_mem_reg[6][7]  ( .D(n2626), .CK(clk), .RN(n4560), .Q(
        \key_mem[6][7] ) );
  DFFRX1 \key_mem_reg[10][7]  ( .D(n3138), .CK(clk), .RN(n4560), .Q(
        \key_mem[10][7] ) );
  DFFRX1 \key_mem_reg[2][6]  ( .D(n2115), .CK(clk), .RN(n4561), .Q(
        \key_mem[2][6] ) );
  DFFRX1 \key_mem_reg[6][6]  ( .D(n2627), .CK(clk), .RN(n4561), .Q(
        \key_mem[6][6] ) );
  DFFRX1 \key_mem_reg[10][6]  ( .D(n3139), .CK(clk), .RN(n4562), .Q(
        \key_mem[10][6] ) );
  DFFRX1 \key_mem_reg[2][5]  ( .D(n2116), .CK(clk), .RN(n4437), .Q(
        \key_mem[2][5] ) );
  DFFRX1 \key_mem_reg[6][5]  ( .D(n2628), .CK(clk), .RN(n4438), .Q(
        \key_mem[6][5] ) );
  DFFRX1 \key_mem_reg[10][5]  ( .D(n3140), .CK(clk), .RN(n4433), .Q(
        \key_mem[10][5] ) );
  DFFRX1 \key_mem_reg[2][4]  ( .D(n2117), .CK(clk), .RN(n4414), .Q(
        \key_mem[2][4] ) );
  DFFRX1 \key_mem_reg[6][4]  ( .D(n2629), .CK(clk), .RN(n4413), .Q(
        \key_mem[6][4] ) );
  DFFRX1 \key_mem_reg[10][4]  ( .D(n3141), .CK(clk), .RN(n4564), .Q(
        \key_mem[10][4] ) );
  DFFRX1 \key_mem_reg[2][3]  ( .D(n2118), .CK(clk), .RN(n4388), .Q(
        \key_mem[2][3] ) );
  DFFRX1 \key_mem_reg[6][3]  ( .D(n2630), .CK(clk), .RN(n4378), .Q(
        \key_mem[6][3] ) );
  DFFRX1 \key_mem_reg[10][3]  ( .D(n3142), .CK(clk), .RN(n4382), .Q(
        \key_mem[10][3] ) );
  DFFRX1 \key_mem_reg[2][2]  ( .D(n2119), .CK(clk), .RN(n4413), .Q(
        \key_mem[2][2] ) );
  DFFRX1 \key_mem_reg[6][2]  ( .D(n2631), .CK(clk), .RN(n4563), .Q(
        \key_mem[6][2] ) );
  DFFRX1 \key_mem_reg[10][2]  ( .D(n3143), .CK(clk), .RN(n4563), .Q(
        \key_mem[10][2] ) );
  DFFRX1 \key_mem_reg[2][1]  ( .D(n2120), .CK(clk), .RN(n4564), .Q(
        \key_mem[2][1] ) );
  DFFRX1 \key_mem_reg[6][1]  ( .D(n2632), .CK(clk), .RN(n4564), .Q(
        \key_mem[6][1] ) );
  DFFRX1 \key_mem_reg[10][1]  ( .D(n3144), .CK(clk), .RN(n4555), .Q(
        \key_mem[10][1] ) );
  DFFRX1 \key_mem_reg[2][0]  ( .D(n2121), .CK(clk), .RN(n4555), .Q(
        \key_mem[2][0] ) );
  DFFRX1 \key_mem_reg[6][0]  ( .D(n2633), .CK(clk), .RN(n4556), .Q(
        \key_mem[6][0] ) );
  DFFRX1 \key_mem_reg[10][0]  ( .D(n3145), .CK(clk), .RN(n4556), .Q(
        \key_mem[10][0] ) );
  DFFRX1 \key_mem_reg[2][127]  ( .D(n1994), .CK(clk), .RN(n4487), .Q(
        \key_mem[2][127] ) );
  DFFRX1 \key_mem_reg[6][127]  ( .D(n2506), .CK(clk), .RN(n4530), .Q(
        \key_mem[6][127] ) );
  DFFRX1 \key_mem_reg[10][127]  ( .D(n3018), .CK(clk), .RN(n4529), .Q(
        \key_mem[10][127] ) );
  DFFRX1 \key_mem_reg[2][95]  ( .D(n2026), .CK(clk), .RN(n4521), .Q(
        \key_mem[2][95] ) );
  DFFRX1 \key_mem_reg[6][95]  ( .D(n2538), .CK(clk), .RN(n4520), .Q(
        \key_mem[6][95] ) );
  DFFRX1 \key_mem_reg[10][95]  ( .D(n3050), .CK(clk), .RN(n4511), .Q(
        \key_mem[10][95] ) );
  DFFRX1 \key_mem_reg[2][63]  ( .D(n2058), .CK(clk), .RN(n4527), .Q(
        \key_mem[2][63] ) );
  DFFRX1 \key_mem_reg[6][63]  ( .D(n2570), .CK(clk), .RN(n4500), .Q(
        \key_mem[6][63] ) );
  DFFRX1 \key_mem_reg[10][63]  ( .D(n3082), .CK(clk), .RN(n4557), .Q(
        \key_mem[10][63] ) );
  DFFRX1 \key_mem_reg[2][31]  ( .D(n2090), .CK(clk), .RN(n4557), .Q(
        \key_mem[2][31] ) );
  DFFRX1 \key_mem_reg[6][31]  ( .D(n2602), .CK(clk), .RN(n4557), .Q(
        \key_mem[6][31] ) );
  DFFRX1 \key_mem_reg[10][31]  ( .D(n3114), .CK(clk), .RN(n4457), .Q(
        \key_mem[10][31] ) );
  DFFRX1 \key_mem_reg[2][120]  ( .D(n2001), .CK(clk), .RN(n4458), .Q(
        \key_mem[2][120] ) );
  DFFRX1 \key_mem_reg[6][120]  ( .D(n2513), .CK(clk), .RN(n4487), .Q(
        \key_mem[6][120] ) );
  DFFRX1 \key_mem_reg[10][120]  ( .D(n3025), .CK(clk), .RN(n4486), .Q(
        \key_mem[10][120] ) );
  DFFRX1 \key_mem_reg[2][88]  ( .D(n2033), .CK(clk), .RN(n4541), .Q(
        \key_mem[2][88] ) );
  DFFRX1 \key_mem_reg[6][88]  ( .D(n2545), .CK(clk), .RN(n4558), .Q(
        \key_mem[6][88] ) );
  DFFRX1 \key_mem_reg[10][88]  ( .D(n3057), .CK(clk), .RN(n4558), .Q(
        \key_mem[10][88] ) );
  DFFRX1 \key_mem_reg[2][56]  ( .D(n2065), .CK(clk), .RN(n4518), .Q(
        \key_mem[2][56] ) );
  DFFRX1 \key_mem_reg[6][56]  ( .D(n2577), .CK(clk), .RN(n4517), .Q(
        \key_mem[6][56] ) );
  DFFRX1 \key_mem_reg[10][56]  ( .D(n3089), .CK(clk), .RN(n4508), .Q(
        \key_mem[10][56] ) );
  DFFRX1 \key_mem_reg[2][24]  ( .D(n2097), .CK(clk), .RN(n4490), .Q(
        \key_mem[2][24] ) );
  DFFRX1 \key_mem_reg[6][24]  ( .D(n2609), .CK(clk), .RN(n4448), .Q(
        \key_mem[6][24] ) );
  DFFRX1 \key_mem_reg[10][24]  ( .D(n3121), .CK(clk), .RN(n4552), .Q(
        \key_mem[10][24] ) );
  DFFRX1 \key_mem_reg[2][122]  ( .D(n1999), .CK(clk), .RN(n4485), .Q(
        \key_mem[2][122] ) );
  DFFRX1 \key_mem_reg[6][122]  ( .D(n2511), .CK(clk), .RN(n4485), .Q(
        \key_mem[6][122] ) );
  DFFRX1 \key_mem_reg[10][122]  ( .D(n3023), .CK(clk), .RN(n4486), .Q(
        \key_mem[10][122] ) );
  DFFRX1 \key_mem_reg[2][90]  ( .D(n2031), .CK(clk), .RN(n4486), .Q(
        \key_mem[2][90] ) );
  DFFRX1 \key_mem_reg[6][90]  ( .D(n2543), .CK(clk), .RN(n4487), .Q(
        \key_mem[6][90] ) );
  DFFRX1 \key_mem_reg[10][90]  ( .D(n3055), .CK(clk), .RN(n4487), .Q(
        \key_mem[10][90] ) );
  DFFRX1 \key_mem_reg[2][58]  ( .D(n2063), .CK(clk), .RN(n4488), .Q(
        \key_mem[2][58] ) );
  DFFRX1 \key_mem_reg[6][58]  ( .D(n2575), .CK(clk), .RN(n4489), .Q(
        \key_mem[6][58] ) );
  DFFRX1 \key_mem_reg[10][58]  ( .D(n3087), .CK(clk), .RN(n4489), .Q(
        \key_mem[10][58] ) );
  DFFRX1 \key_mem_reg[2][26]  ( .D(n2095), .CK(clk), .RN(n4490), .Q(
        \key_mem[2][26] ) );
  DFFRX1 \key_mem_reg[6][26]  ( .D(n2607), .CK(clk), .RN(n4491), .Q(
        \key_mem[6][26] ) );
  DFFRX1 \key_mem_reg[10][26]  ( .D(n3119), .CK(clk), .RN(n4491), .Q(
        \key_mem[10][26] ) );
  DFFRX1 \key_mem_reg[2][123]  ( .D(n1998), .CK(clk), .RN(n4507), .Q(
        \key_mem[2][123] ) );
  DFFRX1 \key_mem_reg[6][123]  ( .D(n2510), .CK(clk), .RN(n4519), .Q(
        \key_mem[6][123] ) );
  DFFRX1 \key_mem_reg[10][123]  ( .D(n3022), .CK(clk), .RN(n4430), .Q(
        \key_mem[10][123] ) );
  DFFRX1 \key_mem_reg[2][91]  ( .D(n2030), .CK(clk), .RN(n4492), .Q(
        \key_mem[2][91] ) );
  DFFRX1 \key_mem_reg[6][91]  ( .D(n2542), .CK(clk), .RN(n4492), .Q(
        \key_mem[6][91] ) );
  DFFRX1 \key_mem_reg[10][91]  ( .D(n3054), .CK(clk), .RN(n4493), .Q(
        \key_mem[10][91] ) );
  DFFRX1 \key_mem_reg[2][59]  ( .D(n2062), .CK(clk), .RN(n4493), .Q(
        \key_mem[2][59] ) );
  DFFRX1 \key_mem_reg[6][59]  ( .D(n2574), .CK(clk), .RN(n4494), .Q(
        \key_mem[6][59] ) );
  DFFRX1 \key_mem_reg[10][59]  ( .D(n3086), .CK(clk), .RN(n4494), .Q(
        \key_mem[10][59] ) );
  DFFRX1 \key_mem_reg[2][27]  ( .D(n2094), .CK(clk), .RN(n4495), .Q(
        \key_mem[2][27] ) );
  DFFRX1 \key_mem_reg[6][27]  ( .D(n2606), .CK(clk), .RN(n4496), .Q(
        \key_mem[6][27] ) );
  DFFRX1 \key_mem_reg[10][27]  ( .D(n3118), .CK(clk), .RN(n4470), .Q(
        \key_mem[10][27] ) );
  DFFRX1 \key_mem_reg[2][126]  ( .D(n1995), .CK(clk), .RN(n4471), .Q(
        \key_mem[2][126] ) );
  DFFRX1 \key_mem_reg[6][126]  ( .D(n2507), .CK(clk), .RN(n4472), .Q(
        \key_mem[6][126] ) );
  DFFRX1 \key_mem_reg[10][126]  ( .D(n3019), .CK(clk), .RN(n4472), .Q(
        \key_mem[10][126] ) );
  DFFRX1 \key_mem_reg[2][94]  ( .D(n2027), .CK(clk), .RN(n4473), .Q(
        \key_mem[2][94] ) );
  DFFRX1 \key_mem_reg[6][94]  ( .D(n2539), .CK(clk), .RN(n4473), .Q(
        \key_mem[6][94] ) );
  DFFRX1 \key_mem_reg[10][94]  ( .D(n3051), .CK(clk), .RN(n4474), .Q(
        \key_mem[10][94] ) );
  DFFRX1 \key_mem_reg[2][62]  ( .D(n2059), .CK(clk), .RN(n4475), .Q(
        \key_mem[2][62] ) );
  DFFRX1 \key_mem_reg[6][62]  ( .D(n2571), .CK(clk), .RN(n4475), .Q(
        \key_mem[6][62] ) );
  DFFRX1 \key_mem_reg[10][62]  ( .D(n3083), .CK(clk), .RN(n4476), .Q(
        \key_mem[10][62] ) );
  DFFRX1 \key_mem_reg[2][30]  ( .D(n2091), .CK(clk), .RN(n4476), .Q(
        \key_mem[2][30] ) );
  DFFRX1 \key_mem_reg[6][30]  ( .D(n2603), .CK(clk), .RN(n4477), .Q(
        \key_mem[6][30] ) );
  DFFRX1 \key_mem_reg[10][30]  ( .D(n3115), .CK(clk), .RN(n4477), .Q(
        \key_mem[10][30] ) );
  DFFRX1 \key_mem_reg[2][125]  ( .D(n1996), .CK(clk), .RN(n4478), .Q(
        \key_mem[2][125] ) );
  DFFRX1 \key_mem_reg[6][125]  ( .D(n2508), .CK(clk), .RN(n4479), .Q(
        \key_mem[6][125] ) );
  DFFRX1 \key_mem_reg[10][125]  ( .D(n3020), .CK(clk), .RN(n4479), .Q(
        \key_mem[10][125] ) );
  DFFRX1 \key_mem_reg[2][93]  ( .D(n2028), .CK(clk), .RN(n4480), .Q(
        \key_mem[2][93] ) );
  DFFRX1 \key_mem_reg[6][93]  ( .D(n2540), .CK(clk), .RN(n4480), .Q(
        \key_mem[6][93] ) );
  DFFRX1 \key_mem_reg[10][93]  ( .D(n3052), .CK(clk), .RN(n4481), .Q(
        \key_mem[10][93] ) );
  DFFRX1 \key_mem_reg[2][61]  ( .D(n2060), .CK(clk), .RN(n4482), .Q(
        \key_mem[2][61] ) );
  DFFRX1 \key_mem_reg[6][61]  ( .D(n2572), .CK(clk), .RN(n4482), .Q(
        \key_mem[6][61] ) );
  DFFRX1 \key_mem_reg[10][61]  ( .D(n3084), .CK(clk), .RN(n4483), .Q(
        \key_mem[10][61] ) );
  DFFRX1 \key_mem_reg[2][29]  ( .D(n2092), .CK(clk), .RN(n4483), .Q(
        \key_mem[2][29] ) );
  DFFRX1 \key_mem_reg[6][29]  ( .D(n2604), .CK(clk), .RN(n4484), .Q(
        \key_mem[6][29] ) );
  DFFRX1 \key_mem_reg[10][29]  ( .D(n3116), .CK(clk), .RN(n4484), .Q(
        \key_mem[10][29] ) );
  DFFRX1 \key_mem_reg[2][124]  ( .D(n1997), .CK(clk), .RN(n4511), .Q(
        \key_mem[2][124] ) );
  DFFRX1 \key_mem_reg[6][124]  ( .D(n2509), .CK(clk), .RN(n4512), .Q(
        \key_mem[6][124] ) );
  DFFRX1 \key_mem_reg[10][124]  ( .D(n3021), .CK(clk), .RN(n4512), .Q(
        \key_mem[10][124] ) );
  DFFRX1 \key_mem_reg[2][92]  ( .D(n2029), .CK(clk), .RN(n4513), .Q(
        \key_mem[2][92] ) );
  DFFRX1 \key_mem_reg[6][92]  ( .D(n2541), .CK(clk), .RN(n4514), .Q(
        \key_mem[6][92] ) );
  DFFRX1 \key_mem_reg[10][92]  ( .D(n3053), .CK(clk), .RN(n4514), .Q(
        \key_mem[10][92] ) );
  DFFRX1 \key_mem_reg[2][60]  ( .D(n2061), .CK(clk), .RN(n4515), .Q(
        \key_mem[2][60] ) );
  DFFRX1 \key_mem_reg[6][60]  ( .D(n2573), .CK(clk), .RN(n4515), .Q(
        \key_mem[6][60] ) );
  DFFRX1 \key_mem_reg[10][60]  ( .D(n3085), .CK(clk), .RN(n4516), .Q(
        \key_mem[10][60] ) );
  DFFRX1 \key_mem_reg[2][28]  ( .D(n2093), .CK(clk), .RN(n4517), .Q(
        \key_mem[2][28] ) );
  DFFRX1 \key_mem_reg[6][28]  ( .D(n2605), .CK(clk), .RN(n4517), .Q(
        \key_mem[6][28] ) );
  DFFRX1 \key_mem_reg[10][28]  ( .D(n3117), .CK(clk), .RN(n4518), .Q(
        \key_mem[10][28] ) );
  DFFRX1 \key_mem_reg[2][121]  ( .D(n2000), .CK(clk), .RN(n4518), .Q(
        \key_mem[2][121] ) );
  DFFRX1 \key_mem_reg[6][121]  ( .D(n2512), .CK(clk), .RN(n4519), .Q(
        \key_mem[6][121] ) );
  DFFRX1 \key_mem_reg[10][121]  ( .D(n3024), .CK(clk), .RN(n4519), .Q(
        \key_mem[10][121] ) );
  DFFRX1 \key_mem_reg[2][89]  ( .D(n2032), .CK(clk), .RN(n4520), .Q(
        \key_mem[2][89] ) );
  DFFRX1 \key_mem_reg[6][89]  ( .D(n2544), .CK(clk), .RN(n4521), .Q(
        \key_mem[6][89] ) );
  DFFRX1 \key_mem_reg[10][89]  ( .D(n3056), .CK(clk), .RN(n4521), .Q(
        \key_mem[10][89] ) );
  DFFRX1 \key_mem_reg[2][57]  ( .D(n2064), .CK(clk), .RN(n4522), .Q(
        \key_mem[2][57] ) );
  DFFRX1 \key_mem_reg[6][57]  ( .D(n2576), .CK(clk), .RN(n4522), .Q(
        \key_mem[6][57] ) );
  DFFRX1 \key_mem_reg[10][57]  ( .D(n3088), .CK(clk), .RN(n4523), .Q(
        \key_mem[10][57] ) );
  DFFRX1 \key_mem_reg[2][25]  ( .D(n2096), .CK(clk), .RN(n4524), .Q(
        \key_mem[2][25] ) );
  DFFRX1 \key_mem_reg[6][25]  ( .D(n2608), .CK(clk), .RN(n4524), .Q(
        \key_mem[6][25] ) );
  DFFRX1 \key_mem_reg[10][25]  ( .D(n3120), .CK(clk), .RN(n4525), .Q(
        \key_mem[10][25] ) );
  DFFRX1 \key_mem_reg[13][119]  ( .D(n3410), .CK(clk), .RN(n4431), .Q(
        \key_mem[13][119] ) );
  DFFRX1 \key_mem_reg[13][118]  ( .D(n3411), .CK(clk), .RN(n4408), .Q(
        \key_mem[13][118] ) );
  DFFRX1 \key_mem_reg[13][117]  ( .D(n3412), .CK(clk), .RN(n4494), .Q(
        \key_mem[13][117] ) );
  DFFRX1 \key_mem_reg[13][116]  ( .D(n3413), .CK(clk), .RN(n4399), .Q(
        \key_mem[13][116] ) );
  DFFRX1 \key_mem_reg[13][115]  ( .D(n3414), .CK(clk), .RN(n4434), .Q(
        \key_mem[13][115] ) );
  DFFRX1 \key_mem_reg[13][114]  ( .D(n3415), .CK(clk), .RN(n4436), .Q(
        \key_mem[13][114] ) );
  DFFRX1 \key_mem_reg[13][113]  ( .D(n3416), .CK(clk), .RN(n4438), .Q(
        \key_mem[13][113] ) );
  DFFRX1 \key_mem_reg[13][112]  ( .D(n3417), .CK(clk), .RN(n4440), .Q(
        \key_mem[13][112] ) );
  DFFRX1 \key_mem_reg[13][111]  ( .D(n3418), .CK(clk), .RN(n4418), .Q(
        \key_mem[13][111] ) );
  DFFRX1 \key_mem_reg[13][110]  ( .D(n3419), .CK(clk), .RN(n4419), .Q(
        \key_mem[13][110] ) );
  DFFRX1 \key_mem_reg[13][109]  ( .D(n3420), .CK(clk), .RN(n4421), .Q(
        \key_mem[13][109] ) );
  DFFRX1 \key_mem_reg[13][108]  ( .D(n3421), .CK(clk), .RN(n4422), .Q(
        \key_mem[13][108] ) );
  DFFRX1 \key_mem_reg[13][106]  ( .D(n3423), .CK(clk), .RN(n4424), .Q(
        \key_mem[13][106] ) );
  DFFRX1 \key_mem_reg[13][105]  ( .D(n3424), .CK(clk), .RN(n4426), .Q(
        \key_mem[13][105] ) );
  DFFRX1 \key_mem_reg[13][104]  ( .D(n3425), .CK(clk), .RN(n4427), .Q(
        \key_mem[13][104] ) );
  DFFRX1 \key_mem_reg[13][103]  ( .D(n3426), .CK(clk), .RN(n4429), .Q(
        \key_mem[13][103] ) );
  DFFRX1 \key_mem_reg[13][102]  ( .D(n3427), .CK(clk), .RN(n4457), .Q(
        \key_mem[13][102] ) );
  DFFRX1 \key_mem_reg[13][101]  ( .D(n3428), .CK(clk), .RN(n4459), .Q(
        \key_mem[13][101] ) );
  DFFRX1 \key_mem_reg[13][100]  ( .D(n3429), .CK(clk), .RN(n4469), .Q(
        \key_mem[13][100] ) );
  DFFRX1 \key_mem_reg[13][99]  ( .D(n3430), .CK(clk), .RN(n4461), .Q(
        \key_mem[13][99] ) );
  DFFRX1 \key_mem_reg[13][98]  ( .D(n3431), .CK(clk), .RN(n4463), .Q(
        \key_mem[13][98] ) );
  DFFRX1 \key_mem_reg[13][97]  ( .D(n3432), .CK(clk), .RN(n4465), .Q(
        \key_mem[13][97] ) );
  DFFRX1 \key_mem_reg[13][96]  ( .D(n3433), .CK(clk), .RN(n4467), .Q(
        \key_mem[13][96] ) );
  DFFRX1 \key_mem_reg[13][87]  ( .D(n3442), .CK(clk), .RN(n4468), .Q(
        \key_mem[13][87] ) );
  DFFRX1 \key_mem_reg[13][86]  ( .D(n3443), .CK(clk), .RN(n4441), .Q(
        \key_mem[13][86] ) );
  DFFRX1 \key_mem_reg[13][85]  ( .D(n3444), .CK(clk), .RN(n4443), .Q(
        \key_mem[13][85] ) );
  DFFRX1 \key_mem_reg[13][84]  ( .D(n3445), .CK(clk), .RN(n4444), .Q(
        \key_mem[13][84] ) );
  DFFRX1 \key_mem_reg[13][83]  ( .D(n3446), .CK(clk), .RN(n4446), .Q(
        \key_mem[13][83] ) );
  DFFRX1 \key_mem_reg[13][82]  ( .D(n3447), .CK(clk), .RN(n4448), .Q(
        \key_mem[13][82] ) );
  DFFRX1 \key_mem_reg[13][81]  ( .D(n3448), .CK(clk), .RN(n4450), .Q(
        \key_mem[13][81] ) );
  DFFRX1 \key_mem_reg[13][80]  ( .D(n3449), .CK(clk), .RN(n4452), .Q(
        \key_mem[13][80] ) );
  DFFRX1 \key_mem_reg[13][79]  ( .D(n3450), .CK(clk), .RN(n4453), .Q(
        \key_mem[13][79] ) );
  DFFRX1 \key_mem_reg[13][78]  ( .D(n3451), .CK(clk), .RN(n4455), .Q(
        \key_mem[13][78] ) );
  DFFRX1 \key_mem_reg[13][77]  ( .D(n3452), .CK(clk), .RN(n4374), .Q(
        \key_mem[13][77] ) );
  DFFRX1 \key_mem_reg[13][76]  ( .D(n3453), .CK(clk), .RN(n4376), .Q(
        \key_mem[13][76] ) );
  DFFRX1 \key_mem_reg[13][75]  ( .D(n3454), .CK(clk), .RN(n4377), .Q(
        \key_mem[13][75] ) );
  DFFRX1 \key_mem_reg[13][74]  ( .D(n3455), .CK(clk), .RN(n4379), .Q(
        \key_mem[13][74] ) );
  DFFRX1 \key_mem_reg[13][73]  ( .D(n3456), .CK(clk), .RN(n4381), .Q(
        \key_mem[13][73] ) );
  DFFRX1 \key_mem_reg[13][72]  ( .D(n3457), .CK(clk), .RN(n4383), .Q(
        \key_mem[13][72] ) );
  DFFRX1 \key_mem_reg[13][71]  ( .D(n3458), .CK(clk), .RN(n4384), .Q(
        \key_mem[13][71] ) );
  DFFRX1 \key_mem_reg[13][70]  ( .D(n3459), .CK(clk), .RN(n4386), .Q(
        \key_mem[13][70] ) );
  DFFRX1 \key_mem_reg[13][69]  ( .D(n3460), .CK(clk), .RN(n4500), .Q(
        \key_mem[13][69] ) );
  DFFRX1 \key_mem_reg[13][68]  ( .D(n3461), .CK(clk), .RN(n4382), .Q(
        \key_mem[13][68] ) );
  DFFRX1 \key_mem_reg[13][67]  ( .D(n3462), .CK(clk), .RN(n4372), .Q(
        \key_mem[13][67] ) );
  DFFRX1 \key_mem_reg[13][66]  ( .D(n3463), .CK(clk), .RN(n4391), .Q(
        \key_mem[13][66] ) );
  DFFRX1 \key_mem_reg[13][65]  ( .D(n3464), .CK(clk), .RN(n4443), .Q(
        \key_mem[13][65] ) );
  DFFRX1 \key_mem_reg[13][64]  ( .D(n3465), .CK(clk), .RN(n4562), .Q(
        \key_mem[13][64] ) );
  DFFRX1 \key_mem_reg[13][55]  ( .D(n3474), .CK(clk), .RN(n4549), .Q(
        \key_mem[13][55] ) );
  DFFRX1 \key_mem_reg[13][54]  ( .D(n3475), .CK(clk), .RN(n4370), .Q(
        \key_mem[13][54] ) );
  DFFRX1 \key_mem_reg[13][53]  ( .D(n3476), .CK(clk), .RN(n4372), .Q(
        \key_mem[13][53] ) );
  DFFRX1 \key_mem_reg[13][52]  ( .D(n3477), .CK(clk), .RN(n4404), .Q(
        \key_mem[13][52] ) );
  DFFRX1 \key_mem_reg[13][51]  ( .D(n3478), .CK(clk), .RN(n4406), .Q(
        \key_mem[13][51] ) );
  DFFRX1 \key_mem_reg[13][50]  ( .D(n3479), .CK(clk), .RN(n4407), .Q(
        \key_mem[13][50] ) );
  DFFRX1 \key_mem_reg[13][49]  ( .D(n3480), .CK(clk), .RN(n4409), .Q(
        \key_mem[13][49] ) );
  DFFRX1 \key_mem_reg[13][47]  ( .D(n3482), .CK(clk), .RN(n4413), .Q(
        \key_mem[13][47] ) );
  DFFRX1 \key_mem_reg[13][46]  ( .D(n3483), .CK(clk), .RN(n4376), .Q(
        \key_mem[13][46] ) );
  DFFRX1 \key_mem_reg[13][45]  ( .D(n3484), .CK(clk), .RN(n4415), .Q(
        \key_mem[13][45] ) );
  DFFRX1 \key_mem_reg[13][44]  ( .D(n3485), .CK(clk), .RN(n4417), .Q(
        \key_mem[13][44] ) );
  DFFRX1 \key_mem_reg[13][43]  ( .D(n3486), .CK(clk), .RN(n4389), .Q(
        \key_mem[13][43] ) );
  DFFRX1 \key_mem_reg[13][42]  ( .D(n3487), .CK(clk), .RN(n4391), .Q(
        \key_mem[13][42] ) );
  DFFRX1 \key_mem_reg[13][41]  ( .D(n3488), .CK(clk), .RN(n4393), .Q(
        \key_mem[13][41] ) );
  DFFRX1 \key_mem_reg[13][40]  ( .D(n3489), .CK(clk), .RN(n4395), .Q(
        \key_mem[13][40] ) );
  DFFRX1 \key_mem_reg[13][39]  ( .D(n3490), .CK(clk), .RN(n4397), .Q(
        \key_mem[13][39] ) );
  DFFRX1 \key_mem_reg[13][38]  ( .D(n3491), .CK(clk), .RN(n4398), .Q(
        \key_mem[13][38] ) );
  DFFRX1 \key_mem_reg[13][37]  ( .D(n3492), .CK(clk), .RN(n4400), .Q(
        \key_mem[13][37] ) );
  DFFRX1 \key_mem_reg[13][36]  ( .D(n3493), .CK(clk), .RN(n4402), .Q(
        \key_mem[13][36] ) );
  DFFRX1 \key_mem_reg[13][35]  ( .D(n3494), .CK(clk), .RN(n4541), .Q(
        \key_mem[13][35] ) );
  DFFRX1 \key_mem_reg[13][34]  ( .D(n3495), .CK(clk), .RN(n4543), .Q(
        \key_mem[13][34] ) );
  DFFRX1 \key_mem_reg[13][33]  ( .D(n3496), .CK(clk), .RN(n4545), .Q(
        \key_mem[13][33] ) );
  DFFRX1 \key_mem_reg[13][32]  ( .D(n3497), .CK(clk), .RN(n4547), .Q(
        \key_mem[13][32] ) );
  DFFRX1 \key_mem_reg[13][23]  ( .D(n3506), .CK(clk), .RN(n4548), .Q(
        \key_mem[13][23] ) );
  DFFRX1 \key_mem_reg[13][22]  ( .D(n3507), .CK(clk), .RN(n4550), .Q(
        \key_mem[13][22] ) );
  DFFRX1 \key_mem_reg[13][21]  ( .D(n3508), .CK(clk), .RN(n4552), .Q(
        \key_mem[13][21] ) );
  DFFRX1 \key_mem_reg[13][20]  ( .D(n3509), .CK(clk), .RN(n4419), .Q(
        \key_mem[13][20] ) );
  DFFRX1 \key_mem_reg[13][18]  ( .D(n3511), .CK(clk), .RN(n4527), .Q(
        \key_mem[13][18] ) );
  DFFRX1 \key_mem_reg[13][16]  ( .D(n3513), .CK(clk), .RN(n4531), .Q(
        \key_mem[13][16] ) );
  DFFRX1 \key_mem_reg[13][15]  ( .D(n3514), .CK(clk), .RN(n4532), .Q(
        \key_mem[13][15] ) );
  DFFRX1 \key_mem_reg[13][14]  ( .D(n3515), .CK(clk), .RN(n4534), .Q(
        \key_mem[13][14] ) );
  DFFRX1 \key_mem_reg[13][13]  ( .D(n3516), .CK(clk), .RN(n4536), .Q(
        \key_mem[13][13] ) );
  DFFRX1 \key_mem_reg[13][12]  ( .D(n3517), .CK(clk), .RN(n4538), .Q(
        \key_mem[13][12] ) );
  DFFRX1 \key_mem_reg[13][11]  ( .D(n3518), .CK(clk), .RN(n4539), .Q(
        \key_mem[13][11] ) );
  DFFRX1 \key_mem_reg[13][10]  ( .D(n3519), .CK(clk), .RN(n4541), .Q(
        \key_mem[13][10] ) );
  DFFRX1 \key_mem_reg[13][9]  ( .D(n3520), .CK(clk), .RN(n4563), .Q(
        \key_mem[13][9] ) );
  DFFRX1 \key_mem_reg[13][8]  ( .D(n3521), .CK(clk), .RN(n4559), .Q(
        \key_mem[13][8] ) );
  DFFRX1 \key_mem_reg[13][7]  ( .D(n3522), .CK(clk), .RN(n4561), .Q(
        \key_mem[13][7] ) );
  DFFRX1 \key_mem_reg[13][6]  ( .D(n3523), .CK(clk), .RN(n4562), .Q(
        \key_mem[13][6] ) );
  DFFRX1 \key_mem_reg[13][5]  ( .D(n3524), .CK(clk), .RN(n4427), .Q(
        \key_mem[13][5] ) );
  DFFRX1 \key_mem_reg[13][4]  ( .D(n3525), .CK(clk), .RN(n4462), .Q(
        \key_mem[13][4] ) );
  DFFRX1 \key_mem_reg[13][3]  ( .D(n3526), .CK(clk), .RN(n4415), .Q(
        \key_mem[13][3] ) );
  DFFRX1 \key_mem_reg[13][2]  ( .D(n3527), .CK(clk), .RN(n4563), .Q(
        \key_mem[13][2] ) );
  DFFRX1 \key_mem_reg[13][1]  ( .D(n3528), .CK(clk), .RN(n4555), .Q(
        \key_mem[13][1] ) );
  DFFRX1 \key_mem_reg[13][0]  ( .D(n3529), .CK(clk), .RN(n4486), .Q(
        \key_mem[13][0] ) );
  DFFRX1 \key_mem_reg[13][127]  ( .D(n3402), .CK(clk), .RN(n4517), .Q(
        \key_mem[13][127] ) );
  DFFRX1 \key_mem_reg[13][95]  ( .D(n3434), .CK(clk), .RN(n4510), .Q(
        \key_mem[13][95] ) );
  DFFRX1 \key_mem_reg[13][63]  ( .D(n3466), .CK(clk), .RN(n4506), .Q(
        \key_mem[13][63] ) );
  DFFRX1 \key_mem_reg[13][31]  ( .D(n3498), .CK(clk), .RN(n4455), .Q(
        \key_mem[13][31] ) );
  DFFRX1 \key_mem_reg[13][120]  ( .D(n3409), .CK(clk), .RN(n4540), .Q(
        \key_mem[13][120] ) );
  DFFRX1 \key_mem_reg[13][88]  ( .D(n3441), .CK(clk), .RN(n4516), .Q(
        \key_mem[13][88] ) );
  DFFRX1 \key_mem_reg[13][56]  ( .D(n3473), .CK(clk), .RN(n4507), .Q(
        \key_mem[13][56] ) );
  DFFRX1 \key_mem_reg[13][24]  ( .D(n3505), .CK(clk), .RN(n4551), .Q(
        \key_mem[13][24] ) );
  DFFRX1 \key_mem_reg[13][122]  ( .D(n3407), .CK(clk), .RN(n4486), .Q(
        \key_mem[13][122] ) );
  DFFRX1 \key_mem_reg[13][90]  ( .D(n3439), .CK(clk), .RN(n4488), .Q(
        \key_mem[13][90] ) );
  DFFRX1 \key_mem_reg[13][58]  ( .D(n3471), .CK(clk), .RN(n4490), .Q(
        \key_mem[13][58] ) );
  DFFRX1 \key_mem_reg[13][26]  ( .D(n3503), .CK(clk), .RN(n4491), .Q(
        \key_mem[13][26] ) );
  DFFRX1 \key_mem_reg[13][123]  ( .D(n3406), .CK(clk), .RN(n4427), .Q(
        \key_mem[13][123] ) );
  DFFRX1 \key_mem_reg[13][91]  ( .D(n3438), .CK(clk), .RN(n4493), .Q(
        \key_mem[13][91] ) );
  DFFRX1 \key_mem_reg[13][59]  ( .D(n3470), .CK(clk), .RN(n4495), .Q(
        \key_mem[13][59] ) );
  DFFRX1 \key_mem_reg[13][27]  ( .D(n3502), .CK(clk), .RN(n4470), .Q(
        \key_mem[13][27] ) );
  DFFRX1 \key_mem_reg[13][126]  ( .D(n3403), .CK(clk), .RN(n4472), .Q(
        \key_mem[13][126] ) );
  DFFRX1 \key_mem_reg[13][94]  ( .D(n3435), .CK(clk), .RN(n4474), .Q(
        \key_mem[13][94] ) );
  DFFRX1 \key_mem_reg[13][62]  ( .D(n3467), .CK(clk), .RN(n4476), .Q(
        \key_mem[13][62] ) );
  DFFRX1 \key_mem_reg[13][30]  ( .D(n3499), .CK(clk), .RN(n4478), .Q(
        \key_mem[13][30] ) );
  DFFRX1 \key_mem_reg[13][125]  ( .D(n3404), .CK(clk), .RN(n4480), .Q(
        \key_mem[13][125] ) );
  DFFRX1 \key_mem_reg[13][93]  ( .D(n3436), .CK(clk), .RN(n4481), .Q(
        \key_mem[13][93] ) );
  DFFRX1 \key_mem_reg[13][61]  ( .D(n3468), .CK(clk), .RN(n4483), .Q(
        \key_mem[13][61] ) );
  DFFRX1 \key_mem_reg[13][29]  ( .D(n3500), .CK(clk), .RN(n4518), .Q(
        \key_mem[13][29] ) );
  DFFRX1 \key_mem_reg[13][124]  ( .D(n3405), .CK(clk), .RN(n4513), .Q(
        \key_mem[13][124] ) );
  DFFRX1 \key_mem_reg[13][92]  ( .D(n3437), .CK(clk), .RN(n4514), .Q(
        \key_mem[13][92] ) );
  DFFRX1 \key_mem_reg[13][60]  ( .D(n3469), .CK(clk), .RN(n4516), .Q(
        \key_mem[13][60] ) );
  DFFRX1 \key_mem_reg[13][28]  ( .D(n3501), .CK(clk), .RN(n4518), .Q(
        \key_mem[13][28] ) );
  DFFRX1 \key_mem_reg[13][121]  ( .D(n3408), .CK(clk), .RN(n4520), .Q(
        \key_mem[13][121] ) );
  DFFRX1 \key_mem_reg[13][89]  ( .D(n3440), .CK(clk), .RN(n4522), .Q(
        \key_mem[13][89] ) );
  DFFRX1 \key_mem_reg[13][57]  ( .D(n3472), .CK(clk), .RN(n4523), .Q(
        \key_mem[13][57] ) );
  DFFRX1 \key_mem_reg[13][25]  ( .D(n3504), .CK(clk), .RN(n4525), .Q(
        \key_mem[13][25] ) );
  DFFRX1 \key_mem_reg[12][119]  ( .D(n3282), .CK(clk), .RN(n4431), .Q(
        \key_mem[12][119] ) );
  DFFRX1 \key_mem_reg[12][118]  ( .D(n3283), .CK(clk), .RN(n4407), .Q(
        \key_mem[12][118] ) );
  DFFRX1 \key_mem_reg[12][117]  ( .D(n3284), .CK(clk), .RN(n4493), .Q(
        \key_mem[12][117] ) );
  DFFRX1 \key_mem_reg[12][116]  ( .D(n3285), .CK(clk), .RN(n4398), .Q(
        \key_mem[12][116] ) );
  DFFRX1 \key_mem_reg[12][115]  ( .D(n3286), .CK(clk), .RN(n4434), .Q(
        \key_mem[12][115] ) );
  DFFRX1 \key_mem_reg[12][114]  ( .D(n3287), .CK(clk), .RN(n4436), .Q(
        \key_mem[12][114] ) );
  DFFRX1 \key_mem_reg[12][113]  ( .D(n3288), .CK(clk), .RN(n4438), .Q(
        \key_mem[12][113] ) );
  DFFRX1 \key_mem_reg[12][112]  ( .D(n3289), .CK(clk), .RN(n4439), .Q(
        \key_mem[12][112] ) );
  DFFRX1 \key_mem_reg[12][111]  ( .D(n3290), .CK(clk), .RN(n4418), .Q(
        \key_mem[12][111] ) );
  DFFRX1 \key_mem_reg[12][110]  ( .D(n3291), .CK(clk), .RN(n4419), .Q(
        \key_mem[12][110] ) );
  DFFRX1 \key_mem_reg[12][109]  ( .D(n3292), .CK(clk), .RN(n4420), .Q(
        \key_mem[12][109] ) );
  DFFRX1 \key_mem_reg[12][108]  ( .D(n3293), .CK(clk), .RN(n4422), .Q(
        \key_mem[12][108] ) );
  DFFRX1 \key_mem_reg[12][106]  ( .D(n3295), .CK(clk), .RN(n4424), .Q(
        \key_mem[12][106] ) );
  DFFRX1 \key_mem_reg[12][105]  ( .D(n3296), .CK(clk), .RN(n4426), .Q(
        \key_mem[12][105] ) );
  DFFRX1 \key_mem_reg[12][104]  ( .D(n3297), .CK(clk), .RN(n4427), .Q(
        \key_mem[12][104] ) );
  DFFRX1 \key_mem_reg[12][103]  ( .D(n3298), .CK(clk), .RN(n4429), .Q(
        \key_mem[12][103] ) );
  DFFRX1 \key_mem_reg[12][102]  ( .D(n3299), .CK(clk), .RN(n4457), .Q(
        \key_mem[12][102] ) );
  DFFRX1 \key_mem_reg[12][101]  ( .D(n3300), .CK(clk), .RN(n4459), .Q(
        \key_mem[12][101] ) );
  DFFRX1 \key_mem_reg[12][100]  ( .D(n3301), .CK(clk), .RN(n4460), .Q(
        \key_mem[12][100] ) );
  DFFRX1 \key_mem_reg[12][99]  ( .D(n3302), .CK(clk), .RN(n4461), .Q(
        \key_mem[12][99] ) );
  DFFRX1 \key_mem_reg[12][98]  ( .D(n3303), .CK(clk), .RN(n4463), .Q(
        \key_mem[12][98] ) );
  DFFRX1 \key_mem_reg[12][97]  ( .D(n3304), .CK(clk), .RN(n4465), .Q(
        \key_mem[12][97] ) );
  DFFRX1 \key_mem_reg[12][96]  ( .D(n3305), .CK(clk), .RN(n4467), .Q(
        \key_mem[12][96] ) );
  DFFRX1 \key_mem_reg[12][87]  ( .D(n3314), .CK(clk), .RN(n4468), .Q(
        \key_mem[12][87] ) );
  DFFRX1 \key_mem_reg[12][86]  ( .D(n3315), .CK(clk), .RN(n4441), .Q(
        \key_mem[12][86] ) );
  DFFRX1 \key_mem_reg[12][85]  ( .D(n3316), .CK(clk), .RN(n4443), .Q(
        \key_mem[12][85] ) );
  DFFRX1 \key_mem_reg[12][84]  ( .D(n3317), .CK(clk), .RN(n4444), .Q(
        \key_mem[12][84] ) );
  DFFRX1 \key_mem_reg[12][83]  ( .D(n3318), .CK(clk), .RN(n4446), .Q(
        \key_mem[12][83] ) );
  DFFRX1 \key_mem_reg[12][82]  ( .D(n3319), .CK(clk), .RN(n4448), .Q(
        \key_mem[12][82] ) );
  DFFRX1 \key_mem_reg[12][81]  ( .D(n3320), .CK(clk), .RN(n4450), .Q(
        \key_mem[12][81] ) );
  DFFRX1 \key_mem_reg[12][80]  ( .D(n3321), .CK(clk), .RN(n4451), .Q(
        \key_mem[12][80] ) );
  DFFRX1 \key_mem_reg[12][79]  ( .D(n3322), .CK(clk), .RN(n4453), .Q(
        \key_mem[12][79] ) );
  DFFRX1 \key_mem_reg[12][78]  ( .D(n3323), .CK(clk), .RN(n4455), .Q(
        \key_mem[12][78] ) );
  DFFRX1 \key_mem_reg[12][77]  ( .D(n3324), .CK(clk), .RN(n4374), .Q(
        \key_mem[12][77] ) );
  DFFRX1 \key_mem_reg[12][76]  ( .D(n3325), .CK(clk), .RN(n4375), .Q(
        \key_mem[12][76] ) );
  DFFRX1 \key_mem_reg[12][75]  ( .D(n3326), .CK(clk), .RN(n4377), .Q(
        \key_mem[12][75] ) );
  DFFRX1 \key_mem_reg[12][74]  ( .D(n3327), .CK(clk), .RN(n4379), .Q(
        \key_mem[12][74] ) );
  DFFRX1 \key_mem_reg[12][73]  ( .D(n3328), .CK(clk), .RN(n4381), .Q(
        \key_mem[12][73] ) );
  DFFRX1 \key_mem_reg[12][72]  ( .D(n3329), .CK(clk), .RN(n4383), .Q(
        \key_mem[12][72] ) );
  DFFRX1 \key_mem_reg[12][71]  ( .D(n3330), .CK(clk), .RN(n4384), .Q(
        \key_mem[12][71] ) );
  DFFRX1 \key_mem_reg[12][70]  ( .D(n3331), .CK(clk), .RN(n4386), .Q(
        \key_mem[12][70] ) );
  DFFRX1 \key_mem_reg[12][69]  ( .D(n3332), .CK(clk), .RN(n4426), .Q(
        \key_mem[12][69] ) );
  DFFRX1 \key_mem_reg[12][68]  ( .D(n3333), .CK(clk), .RN(n4449), .Q(
        \key_mem[12][68] ) );
  DFFRX1 \key_mem_reg[12][67]  ( .D(n3334), .CK(clk), .RN(n4371), .Q(
        \key_mem[12][67] ) );
  DFFRX1 \key_mem_reg[12][66]  ( .D(n3335), .CK(clk), .RN(n4394), .Q(
        \key_mem[12][66] ) );
  DFFRX1 \key_mem_reg[12][65]  ( .D(n3336), .CK(clk), .RN(n4444), .Q(
        \key_mem[12][65] ) );
  DFFRX1 \key_mem_reg[12][64]  ( .D(n3337), .CK(clk), .RN(n4561), .Q(
        \key_mem[12][64] ) );
  DFFRX1 \key_mem_reg[12][55]  ( .D(n3346), .CK(clk), .RN(n4550), .Q(
        \key_mem[12][55] ) );
  DFFRX1 \key_mem_reg[12][54]  ( .D(n3347), .CK(clk), .RN(n4370), .Q(
        \key_mem[12][54] ) );
  DFFRX1 \key_mem_reg[12][53]  ( .D(n3348), .CK(clk), .RN(n4372), .Q(
        \key_mem[12][53] ) );
  DFFRX1 \key_mem_reg[12][52]  ( .D(n3349), .CK(clk), .RN(n4404), .Q(
        \key_mem[12][52] ) );
  DFFRX1 \key_mem_reg[12][51]  ( .D(n3350), .CK(clk), .RN(n4405), .Q(
        \key_mem[12][51] ) );
  DFFRX1 \key_mem_reg[12][50]  ( .D(n3351), .CK(clk), .RN(n4407), .Q(
        \key_mem[12][50] ) );
  DFFRX1 \key_mem_reg[12][49]  ( .D(n3352), .CK(clk), .RN(n4409), .Q(
        \key_mem[12][49] ) );
  DFFRX1 \key_mem_reg[12][47]  ( .D(n3354), .CK(clk), .RN(n4413), .Q(
        \key_mem[12][47] ) );
  DFFRX1 \key_mem_reg[12][46]  ( .D(n3355), .CK(clk), .RN(n4386), .Q(
        \key_mem[12][46] ) );
  DFFRX1 \key_mem_reg[12][45]  ( .D(n3356), .CK(clk), .RN(n4415), .Q(
        \key_mem[12][45] ) );
  DFFRX1 \key_mem_reg[12][44]  ( .D(n3357), .CK(clk), .RN(n4417), .Q(
        \key_mem[12][44] ) );
  DFFRX1 \key_mem_reg[12][43]  ( .D(n3358), .CK(clk), .RN(n4389), .Q(
        \key_mem[12][43] ) );
  DFFRX1 \key_mem_reg[12][42]  ( .D(n3359), .CK(clk), .RN(n4391), .Q(
        \key_mem[12][42] ) );
  DFFRX1 \key_mem_reg[12][41]  ( .D(n3360), .CK(clk), .RN(n4393), .Q(
        \key_mem[12][41] ) );
  DFFRX1 \key_mem_reg[12][40]  ( .D(n3361), .CK(clk), .RN(n4395), .Q(
        \key_mem[12][40] ) );
  DFFRX1 \key_mem_reg[12][39]  ( .D(n3362), .CK(clk), .RN(n4396), .Q(
        \key_mem[12][39] ) );
  DFFRX1 \key_mem_reg[12][38]  ( .D(n3363), .CK(clk), .RN(n4398), .Q(
        \key_mem[12][38] ) );
  DFFRX1 \key_mem_reg[12][37]  ( .D(n3364), .CK(clk), .RN(n4400), .Q(
        \key_mem[12][37] ) );
  DFFRX1 \key_mem_reg[12][36]  ( .D(n3365), .CK(clk), .RN(n4402), .Q(
        \key_mem[12][36] ) );
  DFFRX1 \key_mem_reg[12][35]  ( .D(n3366), .CK(clk), .RN(n4541), .Q(
        \key_mem[12][35] ) );
  DFFRX1 \key_mem_reg[12][34]  ( .D(n3367), .CK(clk), .RN(n4543), .Q(
        \key_mem[12][34] ) );
  DFFRX1 \key_mem_reg[12][33]  ( .D(n3368), .CK(clk), .RN(n4545), .Q(
        \key_mem[12][33] ) );
  DFFRX1 \key_mem_reg[12][32]  ( .D(n3369), .CK(clk), .RN(n4547), .Q(
        \key_mem[12][32] ) );
  DFFRX1 \key_mem_reg[12][23]  ( .D(n3378), .CK(clk), .RN(n4548), .Q(
        \key_mem[12][23] ) );
  DFFRX1 \key_mem_reg[12][22]  ( .D(n3379), .CK(clk), .RN(n4550), .Q(
        \key_mem[12][22] ) );
  DFFRX1 \key_mem_reg[12][21]  ( .D(n3380), .CK(clk), .RN(n4552), .Q(
        \key_mem[12][21] ) );
  DFFRX1 \key_mem_reg[12][20]  ( .D(n3381), .CK(clk), .RN(n4420), .Q(
        \key_mem[12][20] ) );
  DFFRX1 \key_mem_reg[12][18]  ( .D(n3383), .CK(clk), .RN(n4527), .Q(
        \key_mem[12][18] ) );
  DFFRX1 \key_mem_reg[12][17]  ( .D(n3384), .CK(clk), .RN(n4529), .Q(
        \key_mem[12][17] ) );
  DFFRX1 \key_mem_reg[12][16]  ( .D(n3385), .CK(clk), .RN(n4530), .Q(
        \key_mem[12][16] ) );
  DFFRX1 \key_mem_reg[12][15]  ( .D(n3386), .CK(clk), .RN(n4532), .Q(
        \key_mem[12][15] ) );
  DFFRX1 \key_mem_reg[12][14]  ( .D(n3387), .CK(clk), .RN(n4534), .Q(
        \key_mem[12][14] ) );
  DFFRX1 \key_mem_reg[12][13]  ( .D(n3388), .CK(clk), .RN(n4536), .Q(
        \key_mem[12][13] ) );
  DFFRX1 \key_mem_reg[12][12]  ( .D(n3389), .CK(clk), .RN(n4538), .Q(
        \key_mem[12][12] ) );
  DFFRX1 \key_mem_reg[12][11]  ( .D(n3390), .CK(clk), .RN(n4539), .Q(
        \key_mem[12][11] ) );
  DFFRX1 \key_mem_reg[12][10]  ( .D(n3391), .CK(clk), .RN(n4541), .Q(
        \key_mem[12][10] ) );
  DFFRX1 \key_mem_reg[12][9]  ( .D(n3392), .CK(clk), .RN(n4524), .Q(
        \key_mem[12][9] ) );
  DFFRX1 \key_mem_reg[12][8]  ( .D(n3393), .CK(clk), .RN(n4559), .Q(
        \key_mem[12][8] ) );
  DFFRX1 \key_mem_reg[12][7]  ( .D(n3394), .CK(clk), .RN(n4560), .Q(
        \key_mem[12][7] ) );
  DFFRX1 \key_mem_reg[12][6]  ( .D(n3395), .CK(clk), .RN(n4562), .Q(
        \key_mem[12][6] ) );
  DFFRX1 \key_mem_reg[12][5]  ( .D(n3396), .CK(clk), .RN(n4428), .Q(
        \key_mem[12][5] ) );
  DFFRX1 \key_mem_reg[12][4]  ( .D(n3397), .CK(clk), .RN(n4463), .Q(
        \key_mem[12][4] ) );
  DFFRX1 \key_mem_reg[12][3]  ( .D(n3398), .CK(clk), .RN(n4414), .Q(
        \key_mem[12][3] ) );
  DFFRX1 \key_mem_reg[12][2]  ( .D(n3399), .CK(clk), .RN(n4563), .Q(
        \key_mem[12][2] ) );
  DFFRX1 \key_mem_reg[12][1]  ( .D(n3400), .CK(clk), .RN(n4555), .Q(
        \key_mem[12][1] ) );
  DFFRX1 \key_mem_reg[12][0]  ( .D(n3401), .CK(clk), .RN(n4485), .Q(
        \key_mem[12][0] ) );
  DFFRX1 \key_mem_reg[12][127]  ( .D(n3274), .CK(clk), .RN(n4526), .Q(
        \key_mem[12][127] ) );
  DFFRX1 \key_mem_reg[12][95]  ( .D(n3306), .CK(clk), .RN(n4509), .Q(
        \key_mem[12][95] ) );
  DFFRX1 \key_mem_reg[12][63]  ( .D(n3338), .CK(clk), .RN(n4516), .Q(
        \key_mem[12][63] ) );
  DFFRX1 \key_mem_reg[12][31]  ( .D(n3370), .CK(clk), .RN(n4456), .Q(
        \key_mem[12][31] ) );
  DFFRX1 \key_mem_reg[12][120]  ( .D(n3281), .CK(clk), .RN(n4539), .Q(
        \key_mem[12][120] ) );
  DFFRX1 \key_mem_reg[12][88]  ( .D(n3313), .CK(clk), .RN(n4558), .Q(
        \key_mem[12][88] ) );
  DFFRX1 \key_mem_reg[12][56]  ( .D(n3345), .CK(clk), .RN(n4506), .Q(
        \key_mem[12][56] ) );
  DFFRX1 \key_mem_reg[12][24]  ( .D(n3377), .CK(clk), .RN(n4550), .Q(
        \key_mem[12][24] ) );
  DFFRX1 \key_mem_reg[12][122]  ( .D(n3279), .CK(clk), .RN(n4486), .Q(
        \key_mem[12][122] ) );
  DFFRX1 \key_mem_reg[12][90]  ( .D(n3311), .CK(clk), .RN(n4488), .Q(
        \key_mem[12][90] ) );
  DFFRX1 \key_mem_reg[12][58]  ( .D(n3343), .CK(clk), .RN(n4489), .Q(
        \key_mem[12][58] ) );
  DFFRX1 \key_mem_reg[12][26]  ( .D(n3375), .CK(clk), .RN(n4491), .Q(
        \key_mem[12][26] ) );
  DFFRX1 \key_mem_reg[12][123]  ( .D(n3278), .CK(clk), .RN(n4428), .Q(
        \key_mem[12][123] ) );
  DFFRX1 \key_mem_reg[12][91]  ( .D(n3310), .CK(clk), .RN(n4493), .Q(
        \key_mem[12][91] ) );
  DFFRX1 \key_mem_reg[12][59]  ( .D(n3342), .CK(clk), .RN(n4495), .Q(
        \key_mem[12][59] ) );
  DFFRX1 \key_mem_reg[12][27]  ( .D(n3374), .CK(clk), .RN(n4470), .Q(
        \key_mem[12][27] ) );
  DFFRX1 \key_mem_reg[12][126]  ( .D(n3275), .CK(clk), .RN(n4472), .Q(
        \key_mem[12][126] ) );
  DFFRX1 \key_mem_reg[12][94]  ( .D(n3307), .CK(clk), .RN(n4474), .Q(
        \key_mem[12][94] ) );
  DFFRX1 \key_mem_reg[12][62]  ( .D(n3339), .CK(clk), .RN(n4476), .Q(
        \key_mem[12][62] ) );
  DFFRX1 \key_mem_reg[12][30]  ( .D(n3371), .CK(clk), .RN(n4478), .Q(
        \key_mem[12][30] ) );
  DFFRX1 \key_mem_reg[12][125]  ( .D(n3276), .CK(clk), .RN(n4479), .Q(
        \key_mem[12][125] ) );
  DFFRX1 \key_mem_reg[12][93]  ( .D(n3308), .CK(clk), .RN(n4481), .Q(
        \key_mem[12][93] ) );
  DFFRX1 \key_mem_reg[12][61]  ( .D(n3340), .CK(clk), .RN(n4483), .Q(
        \key_mem[12][61] ) );
  DFFRX1 \key_mem_reg[12][29]  ( .D(n3372), .CK(clk), .RN(n4445), .Q(
        \key_mem[12][29] ) );
  DFFRX1 \key_mem_reg[12][124]  ( .D(n3277), .CK(clk), .RN(n4513), .Q(
        \key_mem[12][124] ) );
  DFFRX1 \key_mem_reg[12][92]  ( .D(n3309), .CK(clk), .RN(n4514), .Q(
        \key_mem[12][92] ) );
  DFFRX1 \key_mem_reg[12][60]  ( .D(n3341), .CK(clk), .RN(n4516), .Q(
        \key_mem[12][60] ) );
  DFFRX1 \key_mem_reg[12][28]  ( .D(n3373), .CK(clk), .RN(n4518), .Q(
        \key_mem[12][28] ) );
  DFFRX1 \key_mem_reg[12][121]  ( .D(n3280), .CK(clk), .RN(n4520), .Q(
        \key_mem[12][121] ) );
  DFFRX1 \key_mem_reg[12][89]  ( .D(n3312), .CK(clk), .RN(n4521), .Q(
        \key_mem[12][89] ) );
  DFFRX1 \key_mem_reg[12][57]  ( .D(n3344), .CK(clk), .RN(n4523), .Q(
        \key_mem[12][57] ) );
  DFFRX1 \key_mem_reg[12][25]  ( .D(n3376), .CK(clk), .RN(n4525), .Q(
        \key_mem[12][25] ) );
  DFFRX1 \key_mem_reg[14][119]  ( .D(n3538), .CK(clk), .RN(n4431), .Q(
        \key_mem[14][119] ) );
  DFFRX1 \key_mem_reg[14][118]  ( .D(n3539), .CK(clk), .RN(n4406), .Q(
        \key_mem[14][118] ) );
  DFFRX1 \key_mem_reg[14][117]  ( .D(n3540), .CK(clk), .RN(n4492), .Q(
        \key_mem[14][117] ) );
  DFFRX1 \key_mem_reg[14][116]  ( .D(n3541), .CK(clk), .RN(n4391), .Q(
        \key_mem[14][116] ) );
  DFFRX1 \key_mem_reg[14][115]  ( .D(n3542), .CK(clk), .RN(n4434), .Q(
        \key_mem[14][115] ) );
  DFFRX1 \key_mem_reg[14][114]  ( .D(n3543), .CK(clk), .RN(n4436), .Q(
        \key_mem[14][114] ) );
  DFFRX1 \key_mem_reg[14][113]  ( .D(n3544), .CK(clk), .RN(n4438), .Q(
        \key_mem[14][113] ) );
  DFFRX1 \key_mem_reg[14][112]  ( .D(n3545), .CK(clk), .RN(n4440), .Q(
        \key_mem[14][112] ) );
  DFFRX1 \key_mem_reg[14][111]  ( .D(n3546), .CK(clk), .RN(n4418), .Q(
        \key_mem[14][111] ) );
  DFFRX1 \key_mem_reg[14][110]  ( .D(n3547), .CK(clk), .RN(n4419), .Q(
        \key_mem[14][110] ) );
  DFFRX1 \key_mem_reg[14][109]  ( .D(n3548), .CK(clk), .RN(n4421), .Q(
        \key_mem[14][109] ) );
  DFFRX1 \key_mem_reg[14][108]  ( .D(n3549), .CK(clk), .RN(n4422), .Q(
        \key_mem[14][108] ) );
  DFFRX1 \key_mem_reg[14][107]  ( .D(n3550), .CK(clk), .RN(n4472), .Q(
        \key_mem[14][107] ) );
  DFFRX1 \key_mem_reg[14][106]  ( .D(n3551), .CK(clk), .RN(n4424), .Q(
        \key_mem[14][106] ) );
  DFFRX1 \key_mem_reg[14][105]  ( .D(n3552), .CK(clk), .RN(n4426), .Q(
        \key_mem[14][105] ) );
  DFFRX1 \key_mem_reg[14][104]  ( .D(n3553), .CK(clk), .RN(n4428), .Q(
        \key_mem[14][104] ) );
  DFFRX1 \key_mem_reg[14][103]  ( .D(n3554), .CK(clk), .RN(n4462), .Q(
        \key_mem[14][103] ) );
  DFFRX1 \key_mem_reg[14][102]  ( .D(n3555), .CK(clk), .RN(n4457), .Q(
        \key_mem[14][102] ) );
  DFFRX1 \key_mem_reg[14][101]  ( .D(n3556), .CK(clk), .RN(n4459), .Q(
        \key_mem[14][101] ) );
  DFFRX1 \key_mem_reg[14][100]  ( .D(n3557), .CK(clk), .RN(n4468), .Q(
        \key_mem[14][100] ) );
  DFFRX1 \key_mem_reg[14][99]  ( .D(n3558), .CK(clk), .RN(n4461), .Q(
        \key_mem[14][99] ) );
  DFFRX1 \key_mem_reg[14][98]  ( .D(n3559), .CK(clk), .RN(n4463), .Q(
        \key_mem[14][98] ) );
  DFFRX1 \key_mem_reg[14][97]  ( .D(n3560), .CK(clk), .RN(n4465), .Q(
        \key_mem[14][97] ) );
  DFFRX1 \key_mem_reg[14][96]  ( .D(n3561), .CK(clk), .RN(n4467), .Q(
        \key_mem[14][96] ) );
  DFFRX1 \key_mem_reg[14][87]  ( .D(n3570), .CK(clk), .RN(n4469), .Q(
        \key_mem[14][87] ) );
  DFFRX1 \key_mem_reg[14][86]  ( .D(n3571), .CK(clk), .RN(n4441), .Q(
        \key_mem[14][86] ) );
  DFFRX1 \key_mem_reg[14][85]  ( .D(n3572), .CK(clk), .RN(n4443), .Q(
        \key_mem[14][85] ) );
  DFFRX1 \key_mem_reg[14][84]  ( .D(n3573), .CK(clk), .RN(n4445), .Q(
        \key_mem[14][84] ) );
  DFFRX1 \key_mem_reg[14][83]  ( .D(n3574), .CK(clk), .RN(n4446), .Q(
        \key_mem[14][83] ) );
  DFFRX1 \key_mem_reg[14][82]  ( .D(n3575), .CK(clk), .RN(n4448), .Q(
        \key_mem[14][82] ) );
  DFFRX1 \key_mem_reg[14][81]  ( .D(n3576), .CK(clk), .RN(n4450), .Q(
        \key_mem[14][81] ) );
  DFFRX1 \key_mem_reg[14][80]  ( .D(n3577), .CK(clk), .RN(n4452), .Q(
        \key_mem[14][80] ) );
  DFFRX1 \key_mem_reg[14][79]  ( .D(n3578), .CK(clk), .RN(n4453), .Q(
        \key_mem[14][79] ) );
  DFFRX1 \key_mem_reg[14][78]  ( .D(n3579), .CK(clk), .RN(n4455), .Q(
        \key_mem[14][78] ) );
  DFFRX1 \key_mem_reg[14][77]  ( .D(n3580), .CK(clk), .RN(n4374), .Q(
        \key_mem[14][77] ) );
  DFFRX1 \key_mem_reg[14][76]  ( .D(n3581), .CK(clk), .RN(n4376), .Q(
        \key_mem[14][76] ) );
  DFFRX1 \key_mem_reg[14][75]  ( .D(n3582), .CK(clk), .RN(n4377), .Q(
        \key_mem[14][75] ) );
  DFFRX1 \key_mem_reg[14][74]  ( .D(n3583), .CK(clk), .RN(n4379), .Q(
        \key_mem[14][74] ) );
  DFFRX1 \key_mem_reg[14][73]  ( .D(n3584), .CK(clk), .RN(n4381), .Q(
        \key_mem[14][73] ) );
  DFFRX1 \key_mem_reg[14][72]  ( .D(n3585), .CK(clk), .RN(n4383), .Q(
        \key_mem[14][72] ) );
  DFFRX1 \key_mem_reg[14][71]  ( .D(n3586), .CK(clk), .RN(n4385), .Q(
        \key_mem[14][71] ) );
  DFFRX1 \key_mem_reg[14][70]  ( .D(n3587), .CK(clk), .RN(n4386), .Q(
        \key_mem[14][70] ) );
  DFFRX1 \key_mem_reg[14][69]  ( .D(n3588), .CK(clk), .RN(n4501), .Q(
        \key_mem[14][69] ) );
  DFFRX1 \key_mem_reg[14][68]  ( .D(n3589), .CK(clk), .RN(n4384), .Q(
        \key_mem[14][68] ) );
  DFFRX1 \key_mem_reg[14][67]  ( .D(n3590), .CK(clk), .RN(n4370), .Q(
        \key_mem[14][67] ) );
  DFFRX1 \key_mem_reg[14][66]  ( .D(n3591), .CK(clk), .RN(n4393), .Q(
        \key_mem[14][66] ) );
  DFFRX1 \key_mem_reg[14][65]  ( .D(n3592), .CK(clk), .RN(n4441), .Q(
        \key_mem[14][65] ) );
  DFFRX1 \key_mem_reg[14][64]  ( .D(n3593), .CK(clk), .RN(n4560), .Q(
        \key_mem[14][64] ) );
  DFFRX1 \key_mem_reg[14][55]  ( .D(n3602), .CK(clk), .RN(n4536), .Q(
        \key_mem[14][55] ) );
  DFFRX1 \key_mem_reg[14][54]  ( .D(n3603), .CK(clk), .RN(n4370), .Q(
        \key_mem[14][54] ) );
  DFFRX1 \key_mem_reg[14][53]  ( .D(n3604), .CK(clk), .RN(n4372), .Q(
        \key_mem[14][53] ) );
  DFFRX1 \key_mem_reg[14][52]  ( .D(n3605), .CK(clk), .RN(n4404), .Q(
        \key_mem[14][52] ) );
  DFFRX1 \key_mem_reg[14][51]  ( .D(n3606), .CK(clk), .RN(n4406), .Q(
        \key_mem[14][51] ) );
  DFFRX1 \key_mem_reg[14][50]  ( .D(n3607), .CK(clk), .RN(n4407), .Q(
        \key_mem[14][50] ) );
  DFFRX1 \key_mem_reg[14][49]  ( .D(n3608), .CK(clk), .RN(n4409), .Q(
        \key_mem[14][49] ) );
  DFFRX1 \key_mem_reg[14][47]  ( .D(n3610), .CK(clk), .RN(n4413), .Q(
        \key_mem[14][47] ) );
  DFFRX1 \key_mem_reg[14][46]  ( .D(n3611), .CK(clk), .RN(n4414), .Q(
        \key_mem[14][46] ) );
  DFFRX1 \key_mem_reg[14][45]  ( .D(n3612), .CK(clk), .RN(n4415), .Q(
        \key_mem[14][45] ) );
  DFFRX1 \key_mem_reg[14][44]  ( .D(n3613), .CK(clk), .RN(n4395), .Q(
        \key_mem[14][44] ) );
  DFFRX1 \key_mem_reg[14][43]  ( .D(n3614), .CK(clk), .RN(n4390), .Q(
        \key_mem[14][43] ) );
  DFFRX1 \key_mem_reg[14][42]  ( .D(n3615), .CK(clk), .RN(n4391), .Q(
        \key_mem[14][42] ) );
  DFFRX1 \key_mem_reg[14][41]  ( .D(n3616), .CK(clk), .RN(n4393), .Q(
        \key_mem[14][41] ) );
  DFFRX1 \key_mem_reg[14][40]  ( .D(n3617), .CK(clk), .RN(n4395), .Q(
        \key_mem[14][40] ) );
  DFFRX1 \key_mem_reg[14][39]  ( .D(n3618), .CK(clk), .RN(n4397), .Q(
        \key_mem[14][39] ) );
  DFFRX1 \key_mem_reg[14][38]  ( .D(n3619), .CK(clk), .RN(n4398), .Q(
        \key_mem[14][38] ) );
  DFFRX1 \key_mem_reg[14][37]  ( .D(n3620), .CK(clk), .RN(n4400), .Q(
        \key_mem[14][37] ) );
  DFFRX1 \key_mem_reg[14][36]  ( .D(n3621), .CK(clk), .RN(n4402), .Q(
        \key_mem[14][36] ) );
  DFFRX1 \key_mem_reg[14][35]  ( .D(n3622), .CK(clk), .RN(n4542), .Q(
        \key_mem[14][35] ) );
  DFFRX1 \key_mem_reg[14][34]  ( .D(n3623), .CK(clk), .RN(n4543), .Q(
        \key_mem[14][34] ) );
  DFFRX1 \key_mem_reg[14][33]  ( .D(n3624), .CK(clk), .RN(n4545), .Q(
        \key_mem[14][33] ) );
  DFFRX1 \key_mem_reg[14][32]  ( .D(n3625), .CK(clk), .RN(n4547), .Q(
        \key_mem[14][32] ) );
  DFFRX1 \key_mem_reg[14][23]  ( .D(n3634), .CK(clk), .RN(n4549), .Q(
        \key_mem[14][23] ) );
  DFFRX1 \key_mem_reg[14][22]  ( .D(n3635), .CK(clk), .RN(n4550), .Q(
        \key_mem[14][22] ) );
  DFFRX1 \key_mem_reg[14][21]  ( .D(n3636), .CK(clk), .RN(n4552), .Q(
        \key_mem[14][21] ) );
  DFFRX1 \key_mem_reg[14][20]  ( .D(n3637), .CK(clk), .RN(n4418), .Q(
        \key_mem[14][20] ) );
  DFFRX1 \key_mem_reg[14][19]  ( .D(n3638), .CK(clk), .RN(n4554), .Q(
        \key_mem[14][19] ) );
  DFFRX1 \key_mem_reg[14][18]  ( .D(n3639), .CK(clk), .RN(n4527), .Q(
        \key_mem[14][18] ) );
  DFFRX1 \key_mem_reg[14][17]  ( .D(n3640), .CK(clk), .RN(n4529), .Q(
        \key_mem[14][17] ) );
  DFFRX1 \key_mem_reg[14][16]  ( .D(n3641), .CK(clk), .RN(n4531), .Q(
        \key_mem[14][16] ) );
  DFFRX1 \key_mem_reg[14][15]  ( .D(n3642), .CK(clk), .RN(n4532), .Q(
        \key_mem[14][15] ) );
  DFFRX1 \key_mem_reg[14][14]  ( .D(n3643), .CK(clk), .RN(n4534), .Q(
        \key_mem[14][14] ) );
  DFFRX1 \key_mem_reg[14][13]  ( .D(n3644), .CK(clk), .RN(n4536), .Q(
        \key_mem[14][13] ) );
  DFFRX1 \key_mem_reg[14][12]  ( .D(n3645), .CK(clk), .RN(n4538), .Q(
        \key_mem[14][12] ) );
  DFFRX1 \key_mem_reg[14][11]  ( .D(n3646), .CK(clk), .RN(n4540), .Q(
        \key_mem[14][11] ) );
  DFFRX1 \key_mem_reg[14][10]  ( .D(n3647), .CK(clk), .RN(n4439), .Q(
        \key_mem[14][10] ) );
  DFFRX1 \key_mem_reg[14][9]  ( .D(n3648), .CK(clk), .RN(n4525), .Q(
        \key_mem[14][9] ) );
  DFFRX1 \key_mem_reg[14][8]  ( .D(n3649), .CK(clk), .RN(n4559), .Q(
        \key_mem[14][8] ) );
  DFFRX1 \key_mem_reg[14][7]  ( .D(n3650), .CK(clk), .RN(n4561), .Q(
        \key_mem[14][7] ) );
  DFFRX1 \key_mem_reg[14][6]  ( .D(n3651), .CK(clk), .RN(n4562), .Q(
        \key_mem[14][6] ) );
  DFFRX1 \key_mem_reg[14][5]  ( .D(n3652), .CK(clk), .RN(n4430), .Q(
        \key_mem[14][5] ) );
  DFFRX1 \key_mem_reg[14][4]  ( .D(n3653), .CK(clk), .RN(n4465), .Q(
        \key_mem[14][4] ) );
  DFFRX1 \key_mem_reg[14][3]  ( .D(n3654), .CK(clk), .RN(n4416), .Q(
        \key_mem[14][3] ) );
  DFFRX1 \key_mem_reg[14][2]  ( .D(n3655), .CK(clk), .RN(n4564), .Q(
        \key_mem[14][2] ) );
  DFFRX1 \key_mem_reg[14][1]  ( .D(n3656), .CK(clk), .RN(n4555), .Q(
        \key_mem[14][1] ) );
  DFFRX1 \key_mem_reg[14][0]  ( .D(n3657), .CK(clk), .RN(n4484), .Q(
        \key_mem[14][0] ) );
  DFFRX1 \key_mem_reg[14][127]  ( .D(n3530), .CK(clk), .RN(n4518), .Q(
        \key_mem[14][127] ) );
  DFFRX1 \key_mem_reg[14][95]  ( .D(n3562), .CK(clk), .RN(n4508), .Q(
        \key_mem[14][95] ) );
  DFFRX1 \key_mem_reg[14][63]  ( .D(n3594), .CK(clk), .RN(n4525), .Q(
        \key_mem[14][63] ) );
  DFFRX1 \key_mem_reg[14][31]  ( .D(n3626), .CK(clk), .RN(n4453), .Q(
        \key_mem[14][31] ) );
  DFFRX1 \key_mem_reg[14][120]  ( .D(n3537), .CK(clk), .RN(n4556), .Q(
        \key_mem[14][120] ) );
  DFFRX1 \key_mem_reg[14][88]  ( .D(n3569), .CK(clk), .RN(n4515), .Q(
        \key_mem[14][88] ) );
  DFFRX1 \key_mem_reg[14][56]  ( .D(n3601), .CK(clk), .RN(n4505), .Q(
        \key_mem[14][56] ) );
  DFFRX1 \key_mem_reg[14][24]  ( .D(n3633), .CK(clk), .RN(n4549), .Q(
        \key_mem[14][24] ) );
  DFFRX1 \key_mem_reg[14][122]  ( .D(n3535), .CK(clk), .RN(n4486), .Q(
        \key_mem[14][122] ) );
  DFFRX1 \key_mem_reg[14][90]  ( .D(n3567), .CK(clk), .RN(n4488), .Q(
        \key_mem[14][90] ) );
  DFFRX1 \key_mem_reg[14][58]  ( .D(n3599), .CK(clk), .RN(n4490), .Q(
        \key_mem[14][58] ) );
  DFFRX1 \key_mem_reg[14][26]  ( .D(n3631), .CK(clk), .RN(n4528), .Q(
        \key_mem[14][26] ) );
  DFFRX1 \key_mem_reg[14][123]  ( .D(n3534), .CK(clk), .RN(n4425), .Q(
        \key_mem[14][123] ) );
  DFFRX1 \key_mem_reg[14][91]  ( .D(n3566), .CK(clk), .RN(n4493), .Q(
        \key_mem[14][91] ) );
  DFFRX1 \key_mem_reg[14][59]  ( .D(n3598), .CK(clk), .RN(n4495), .Q(
        \key_mem[14][59] ) );
  DFFRX1 \key_mem_reg[14][27]  ( .D(n3630), .CK(clk), .RN(n4470), .Q(
        \key_mem[14][27] ) );
  DFFRX1 \key_mem_reg[14][126]  ( .D(n3531), .CK(clk), .RN(n4473), .Q(
        \key_mem[14][126] ) );
  DFFRX1 \key_mem_reg[14][94]  ( .D(n3563), .CK(clk), .RN(n4474), .Q(
        \key_mem[14][94] ) );
  DFFRX1 \key_mem_reg[14][62]  ( .D(n3595), .CK(clk), .RN(n4476), .Q(
        \key_mem[14][62] ) );
  DFFRX1 \key_mem_reg[14][30]  ( .D(n3627), .CK(clk), .RN(n4478), .Q(
        \key_mem[14][30] ) );
  DFFRX1 \key_mem_reg[14][125]  ( .D(n3532), .CK(clk), .RN(n4480), .Q(
        \key_mem[14][125] ) );
  DFFRX1 \key_mem_reg[14][93]  ( .D(n3564), .CK(clk), .RN(n4481), .Q(
        \key_mem[14][93] ) );
  DFFRX1 \key_mem_reg[14][61]  ( .D(n3596), .CK(clk), .RN(n4483), .Q(
        \key_mem[14][61] ) );
  DFFRX1 \key_mem_reg[14][29]  ( .D(n3628), .CK(clk), .RN(n4511), .Q(
        \key_mem[14][29] ) );
  DFFRX1 \key_mem_reg[14][124]  ( .D(n3533), .CK(clk), .RN(n4513), .Q(
        \key_mem[14][124] ) );
  DFFRX1 \key_mem_reg[14][92]  ( .D(n3565), .CK(clk), .RN(n4515), .Q(
        \key_mem[14][92] ) );
  DFFRX1 \key_mem_reg[14][60]  ( .D(n3597), .CK(clk), .RN(n4516), .Q(
        \key_mem[14][60] ) );
  DFFRX1 \key_mem_reg[14][28]  ( .D(n3629), .CK(clk), .RN(n4518), .Q(
        \key_mem[14][28] ) );
  DFFRX1 \key_mem_reg[14][121]  ( .D(n3536), .CK(clk), .RN(n4520), .Q(
        \key_mem[14][121] ) );
  DFFRX1 \key_mem_reg[14][89]  ( .D(n3568), .CK(clk), .RN(n4522), .Q(
        \key_mem[14][89] ) );
  DFFRX1 \key_mem_reg[14][57]  ( .D(n3600), .CK(clk), .RN(n4523), .Q(
        \key_mem[14][57] ) );
  DFFRX1 \key_mem_reg[14][25]  ( .D(n3632), .CK(clk), .RN(n4525), .Q(
        \key_mem[14][25] ) );
  DFFRX1 \key_mem_reg[12][48]  ( .D(n3353), .CK(clk), .RN(n4411), .Q(
        \key_mem[12][48] ) );
  DFFRX1 \key_mem_reg[1][48]  ( .D(n1945), .CK(clk), .RN(n4505), .Q(
        \key_mem[1][48] ) );
  DFFRX1 \key_mem_reg[5][48]  ( .D(n2457), .CK(clk), .RN(n4410), .Q(
        \key_mem[5][48] ) );
  DFFRX1 \key_mem_reg[9][48]  ( .D(n2969), .CK(clk), .RN(n4410), .Q(
        \key_mem[9][48] ) );
  DFFRX1 \key_mem_reg[13][48]  ( .D(n3481), .CK(clk), .RN(n4411), .Q(
        \key_mem[13][48] ) );
  DFFRX1 \key_mem_reg[8][48]  ( .D(n2841), .CK(clk), .RN(n4410), .Q(
        \key_mem[8][48] ) );
  DFFRX1 \key_mem_reg[4][48]  ( .D(n2329), .CK(clk), .RN(n4410), .Q(
        \key_mem[4][48] ) );
  DFFRX1 \key_mem_reg[0][48]  ( .D(n1817), .CK(clk), .RN(n4409), .Q(
        \key_mem[0][48] ) );
  DFFRX1 \key_mem_reg[10][48]  ( .D(n3097), .CK(clk), .RN(n4411), .Q(
        \key_mem[10][48] ) );
  DFFRX1 \key_mem_reg[6][48]  ( .D(n2585), .CK(clk), .RN(n4410), .Q(
        \key_mem[6][48] ) );
  DFFRX1 \key_mem_reg[2][48]  ( .D(n2073), .CK(clk), .RN(n4409), .Q(
        \key_mem[2][48] ) );
  DFFRX1 \key_mem_reg[11][48]  ( .D(n3225), .CK(clk), .RN(n4411), .Q(
        \key_mem[11][48] ) );
  DFFRX1 \key_mem_reg[3][48]  ( .D(n2201), .CK(clk), .RN(n4410), .Q(
        \key_mem[3][48] ) );
  DFFRX1 \key_mem_reg[7][48]  ( .D(n2713), .CK(clk), .RN(n4410), .Q(
        \key_mem[7][48] ) );
  DFFRX1 \key_mem_reg[9][17]  ( .D(n3000), .CK(clk), .RN(n4528), .Q(
        \key_mem[9][17] ) );
  DFFRX1 \key_mem_reg[5][17]  ( .D(n2488), .CK(clk), .RN(n4528), .Q(
        \key_mem[5][17] ) );
  DFFRX1 \key_mem_reg[11][17]  ( .D(n3256), .CK(clk), .RN(n4529), .Q(
        \key_mem[11][17] ) );
  DFFRX1 \key_mem_reg[7][17]  ( .D(n2744), .CK(clk), .RN(n4528), .Q(
        \key_mem[7][17] ) );
  DFFRX1 \key_mem_reg[3][17]  ( .D(n2232), .CK(clk), .RN(n4528), .Q(
        \key_mem[3][17] ) );
  DFFRX1 \key_mem_reg[13][17]  ( .D(n3512), .CK(clk), .RN(n4529), .Q(
        \key_mem[13][17] ) );
  DFFRX1 \key_mem_reg[14][48]  ( .D(n3609), .CK(clk), .RN(n4411), .Q(
        \key_mem[14][48] ) );
  DFFRX1 \key_mem_ctrl_reg_reg[0]  ( .D(n3927), .CK(clk), .RN(n4470), .Q(
        key_mem_ctrl_reg[0]), .QN(n299) );
  DFFQX1 \prev_key1_reg_reg[31]  ( .D(n3881), .CK(clk), .Q(sboxw[31]) );
  DFFQX1 \prev_key1_reg_reg[30]  ( .D(n3882), .CK(clk), .Q(sboxw[30]) );
  DFFQX1 \prev_key1_reg_reg[23]  ( .D(n3889), .CK(clk), .Q(sboxw[23]) );
  DFFQX1 \prev_key1_reg_reg[22]  ( .D(n3890), .CK(clk), .Q(sboxw[22]) );
  DFFRX1 \key_mem_ctrl_reg_reg[1]  ( .D(n3926), .CK(clk), .RN(n4390), .Q(
        key_mem_ctrl_reg[1]), .QN(n298) );
  DFFRX1 \round_ctr_reg_reg[0]  ( .D(n3925), .CK(clk), .RN(n4429), .Q(
        round_ctr_reg[0]), .QN(n279) );
  DFFQX1 \prev_key1_reg_reg[26]  ( .D(n3886), .CK(clk), .Q(sboxw[26]) );
  DFFQX1 \prev_key1_reg_reg[29]  ( .D(n3883), .CK(clk), .Q(sboxw[29]) );
  DFFQX1 \prev_key1_reg_reg[28]  ( .D(n3884), .CK(clk), .Q(sboxw[28]) );
  DFFQX1 \prev_key1_reg_reg[21]  ( .D(n3891), .CK(clk), .Q(sboxw[21]) );
  DFFQX1 \prev_key1_reg_reg[20]  ( .D(n3892), .CK(clk), .Q(sboxw[20]) );
  DFFQX1 \prev_key1_reg_reg[19]  ( .D(n3893), .CK(clk), .Q(sboxw[19]) );
  DFFQX1 \prev_key1_reg_reg[18]  ( .D(n3894), .CK(clk), .Q(sboxw[18]) );
  DFFQX1 \prev_key1_reg_reg[16]  ( .D(n3896), .CK(clk), .Q(sboxw[16]) );
  DFFQX1 \prev_key1_reg_reg[24]  ( .D(n3888), .CK(clk), .Q(sboxw[24]) );
  DFFQX1 \prev_key1_reg_reg[27]  ( .D(n3885), .CK(clk), .Q(sboxw[27]) );
  DFFQX1 \prev_key1_reg_reg[25]  ( .D(n3887), .CK(clk), .Q(sboxw[25]) );
  DFFQX1 \prev_key1_reg_reg[17]  ( .D(n3895), .CK(clk), .Q(sboxw[17]) );
  DFFQX1 \prev_key1_reg_reg[7]  ( .D(n3905), .CK(clk), .Q(sboxw[7]) );
  DFFQX1 \prev_key1_reg_reg[4]  ( .D(n3908), .CK(clk), .Q(sboxw[4]) );
  DFFQX1 \prev_key1_reg_reg[6]  ( .D(n3906), .CK(clk), .Q(sboxw[6]) );
  DFFQX1 \prev_key1_reg_reg[5]  ( .D(n3907), .CK(clk), .Q(sboxw[5]) );
  DFFQX1 \prev_key1_reg_reg[3]  ( .D(n3909), .CK(clk), .Q(sboxw[3]) );
  DFFQX1 \prev_key1_reg_reg[2]  ( .D(n3910), .CK(clk), .Q(sboxw[2]) );
  DFFQX1 \prev_key1_reg_reg[0]  ( .D(n3912), .CK(clk), .Q(sboxw[0]) );
  DFFQX1 \prev_key1_reg_reg[1]  ( .D(n3911), .CK(clk), .Q(sboxw[1]) );
  DFFQX1 \prev_key1_reg_reg[15]  ( .D(n3897), .CK(clk), .Q(sboxw[15]) );
  DFFQX1 \prev_key1_reg_reg[14]  ( .D(n3898), .CK(clk), .Q(sboxw[14]) );
  DFFQX1 \prev_key1_reg_reg[12]  ( .D(n3900), .CK(clk), .Q(sboxw[12]) );
  DFFQX1 \prev_key1_reg_reg[8]  ( .D(n3904), .CK(clk), .Q(sboxw[8]) );
  DFFQX1 \prev_key1_reg_reg[13]  ( .D(n3899), .CK(clk), .Q(sboxw[13]) );
  DFFQX1 \prev_key1_reg_reg[11]  ( .D(n3901), .CK(clk), .Q(sboxw[11]) );
  DFFQX1 \prev_key1_reg_reg[10]  ( .D(n3902), .CK(clk), .Q(sboxw[10]) );
  DFFQX1 \prev_key1_reg_reg[9]  ( .D(n3903), .CK(clk), .Q(sboxw[9]) );
  DFFRX1 \round_ctr_reg_reg[2]  ( .D(n3923), .CK(clk), .RN(n4429), .Q(
        round_ctr_reg[2]), .QN(n277) );
  DFFRX1 \round_ctr_reg_reg[3]  ( .D(n3922), .CK(clk), .RN(n4430), .Q(
        round_ctr_reg[3]), .QN(n276) );
  DFFRX1 \round_ctr_reg_reg[1]  ( .D(n3924), .CK(clk), .RN(n4440), .Q(
        round_ctr_reg[1]), .QN(n278) );
  OAI221XL U4 ( .A0(n825), .A1(n3998), .B0(n3945), .B1(n5815), .C0(n826), .Y(
        n613) );
  XOR2XL U5 ( .A(n4963), .B(new_sboxw[11]), .Y(n825) );
  XOR2XL U6 ( .A(n4971), .B(new_sboxw[11]), .Y(n4972) );
  XOR2XL U7 ( .A(n4982), .B(new_sboxw[11]), .Y(n4964) );
  XOR2XL U8 ( .A(n4983), .B(new_sboxw[11]), .Y(n4984) );
  INVXL U9 ( .A(new_sboxw[9]), .Y(n5154) );
  XOR2XL U10 ( .A(n5246), .B(new_sboxw[11]), .Y(n5698) );
  XOR2XL U11 ( .A(n5234), .B(new_sboxw[11]), .Y(n5699) );
  XOR2XL U12 ( .A(n5245), .B(new_sboxw[11]), .Y(n5700) );
  XOR2XL U13 ( .A(n4609), .B(new_sboxw[0]), .Y(n869) );
  XOR2XL U14 ( .A(n4883), .B(new_sboxw[0]), .Y(n5732) );
  XNOR2XL U15 ( .A(n5080), .B(new_sboxw[6]), .Y(n4) );
  XNOR2XL U16 ( .A(n4617), .B(new_sboxw[0]), .Y(n3) );
  XOR2XL U17 ( .A(n4627), .B(new_sboxw[0]), .Y(n4610) );
  XOR2XL U18 ( .A(n4897), .B(new_sboxw[9]), .Y(n833) );
  XOR2XL U19 ( .A(n4672), .B(new_sboxw[2]), .Y(n861) );
  XOR2XL U20 ( .A(n4704), .B(new_sboxw[3]), .Y(n857) );
  XOR2XL U21 ( .A(n4768), .B(new_sboxw[5]), .Y(n849) );
  XOR2XL U22 ( .A(n4831), .B(new_sboxw[7]), .Y(n841) );
  XOR2XL U23 ( .A(n4930), .B(new_sboxw[10]), .Y(n829) );
  XOR2XL U24 ( .A(n5029), .B(new_sboxw[13]), .Y(n817) );
  XOR2XL U25 ( .A(n5094), .B(new_sboxw[15]), .Y(n809) );
  XOR2XL U26 ( .A(n5279), .B(new_sboxw[12]), .Y(n5695) );
  XOR2XL U27 ( .A(n5344), .B(new_sboxw[14]), .Y(n5690) );
  XOR2XL U28 ( .A(n5168), .B(new_sboxw[9]), .Y(n5705) );
  XOR2XL U29 ( .A(n4917), .B(new_sboxw[1]), .Y(n5727) );
  XOR2XL U30 ( .A(n4996), .B(new_sboxw[12]), .Y(n821) );
  XOR2XL U31 ( .A(n5062), .B(new_sboxw[14]), .Y(n813) );
  XOR2XL U32 ( .A(n4640), .B(new_sboxw[1]), .Y(n865) );
  XNOR2XL U33 ( .A(n5333), .B(new_sboxw[14]), .Y(n5) );
  XOR2XL U34 ( .A(n4755), .B(new_sboxw[4]), .Y(n4737) );
  XOR2XL U35 ( .A(n5016), .B(new_sboxw[12]), .Y(n5017) );
  XOR2XL U36 ( .A(n5004), .B(new_sboxw[12]), .Y(n5005) );
  XOR2XL U37 ( .A(n5015), .B(new_sboxw[12]), .Y(n4997) );
  XOR2XL U38 ( .A(n5080), .B(new_sboxw[14]), .Y(n5063) );
  XOR2XL U39 ( .A(n4756), .B(new_sboxw[4]), .Y(n4757) );
  XOR2XL U40 ( .A(n4884), .B(new_sboxw[8]), .Y(n4885) );
  XOR2XL U41 ( .A(n4872), .B(new_sboxw[8]), .Y(n4873) );
  AOI222XL U42 ( .A0(n1712), .A1(n7), .B0(key[19]), .B1(n1687), .C0(n1702), 
        .C1(n5698), .Y(n1178) );
  AOI222XL U43 ( .A0(n1710), .A1(n1051), .B0(key[51]), .B1(n1683), .C0(n1697), 
        .C1(n5699), .Y(n1050) );
  AOI222XL U44 ( .A0(n1707), .A1(n6), .B0(key[83]), .B1(n1682), .C0(n5758), 
        .C1(n5700), .Y(n922) );
  NAND2BXL U45 ( .AN(n5762), .B(keylen), .Y(n5678) );
  NAND2BXL U46 ( .AN(n3934), .B(keylen), .Y(n4589) );
  NAND2BXL U47 ( .AN(keylen), .B(n4597), .Y(n4598) );
  XNOR2XL U48 ( .A(round_ctr_reg[2]), .B(keylen), .Y(n75) );
  NAND2BX1 U49 ( .AN(n4565), .B(n1691), .Y(n5674) );
  INVX1 U50 ( .A(n4603), .Y(n5668) );
  NAND2BX1 U51 ( .AN(n4602), .B(n4545), .Y(n5669) );
  INVX1 U52 ( .A(n4599), .Y(n5672) );
  INVX1 U53 ( .A(n4593), .Y(n5758) );
  INVXL U54 ( .A(n5233), .Y(n795) );
  INVXL U55 ( .A(n5244), .Y(n1051) );
  OR2X1 U56 ( .A(n4565), .B(n4589), .Y(n5663) );
  INVX1 U57 ( .A(n4601), .Y(n5671) );
  AOI21X1 U58 ( .A0(n4589), .A1(n4591), .B0(n4565), .Y(n1) );
  INVX1 U59 ( .A(n5678), .Y(n5757) );
  NAND2BX1 U60 ( .AN(n279), .B(n4592), .Y(n742) );
  INVX1 U61 ( .A(n4598), .Y(n5759) );
  OAI221XL U62 ( .A0(n1221), .A1(n3992), .B0(n3935), .B1(n5789), .C0(n1222), 
        .Y(n712) );
  OAI221XL U63 ( .A0(n1197), .A1(n4002), .B0(n3936), .B1(n5869), .C0(n1198), 
        .Y(n706) );
  OAI221XL U64 ( .A0(n869), .A1(n3997), .B0(n3944), .B1(n5796), .C0(n870), .Y(
        n624) );
  OAI221XL U65 ( .A0(n3), .A1(n4003), .B0(n3938), .B1(n5792), .C0(n1126), .Y(
        n688) );
  OAI221XL U66 ( .A0(n1101), .A1(n4000), .B0(n3938), .B1(n5872), .C0(n1102), 
        .Y(n682) );
  OAI221XL U67 ( .A0(n813), .A1(n3999), .B0(n3946), .B1(n5863), .C0(n814), .Y(
        n610) );
  OAI221XL U68 ( .A0(n793), .A1(n3999), .B0(n3946), .B1(n5829), .C0(n794), .Y(
        n605) );
  OAI221XL U69 ( .A0(n837), .A1(n3998), .B0(n3945), .B1(n5783), .C0(n838), .Y(
        n616) );
  OAI221XL U70 ( .A0(n1229), .A1(n3992), .B0(n3935), .B1(n5870), .C0(n1230), 
        .Y(n714) );
  OAI221XL U71 ( .A0(n1049), .A1(n3993), .B0(n3940), .B1(n5825), .C0(n1050), 
        .Y(n669) );
  OAI221XL U72 ( .A0(n921), .A1(n3996), .B0(n3943), .B1(n5827), .C0(n922), .Y(
        n637) );
  OAI221XL U73 ( .A0(n1177), .A1(n4005), .B0(n3936), .B1(n5823), .C0(n1178), 
        .Y(n701) );
  OAI221XL U74 ( .A0(n1209), .A1(n4004), .B0(n3936), .B1(n5821), .C0(n1210), 
        .Y(n709) );
  OAI221XL U75 ( .A0(n973), .A1(n3995), .B0(n3942), .B1(n5874), .C0(n974), .Y(
        n650) );
  OAI221XL U76 ( .A0(n953), .A1(n3995), .B0(n3942), .B1(n5817), .C0(n954), .Y(
        n645) );
  OAI221XL U77 ( .A0(n1081), .A1(n4004), .B0(n3939), .B1(n5819), .C0(n1082), 
        .Y(n677) );
  INVXL U78 ( .A(n5698), .Y(n5250) );
  INVXL U79 ( .A(n5699), .Y(n5238) );
  INVXL U80 ( .A(n5700), .Y(n5230) );
  XOR2XL U81 ( .A(n5220), .B(prev_key0_reg[115]), .Y(n5224) );
  OAI221XL U82 ( .A0(n997), .A1(n3994), .B0(n3941), .B1(n5794), .C0(n998), .Y(
        n656) );
  XNOR2XL U83 ( .A(n5233), .B(prev_key1_reg[83]), .Y(n6) );
  OAI221XL U84 ( .A0(n845), .A1(n3998), .B0(n3945), .B1(n5876), .C0(n846), .Y(
        n618) );
  OAI221XL U85 ( .A0(n1422), .A1(n3992), .B0(n3935), .B1(n5790), .C0(n1254), 
        .Y(n720) );
  OAI221XL U86 ( .A0(n1213), .A1(n4001), .B0(n3936), .B1(n5805), .C0(n1214), 
        .Y(n710) );
  OAI221XL U87 ( .A0(n1201), .A1(n4003), .B0(n3936), .B1(n5853), .C0(n1202), 
        .Y(n707) );
  OAI221XL U88 ( .A0(n1193), .A1(n4004), .B0(n3936), .B1(n5885), .C0(n1194), 
        .Y(n705) );
  OAI221XL U89 ( .A0(n1181), .A1(n4002), .B0(n3936), .B1(n5807), .C0(n1182), 
        .Y(n702) );
  OAI221XL U90 ( .A0(n1169), .A1(n4001), .B0(n3937), .B1(n5855), .C0(n1170), 
        .Y(n699) );
  OAI221XL U91 ( .A0(n1161), .A1(n742), .B0(n3937), .B1(n5887), .C0(n1162), 
        .Y(n697) );
  OAI221XL U92 ( .A0(n1085), .A1(n4003), .B0(n3939), .B1(n5803), .C0(n1086), 
        .Y(n678) );
  OAI221XL U93 ( .A0(n1073), .A1(n742), .B0(n3939), .B1(n5851), .C0(n1074), 
        .Y(n675) );
  OAI221XL U94 ( .A0(n1065), .A1(n4002), .B0(n3939), .B1(n5883), .C0(n1066), 
        .Y(n673) );
  OAI221XL U95 ( .A0(n1053), .A1(n3993), .B0(n3940), .B1(n5809), .C0(n1054), 
        .Y(n670) );
  OAI221XL U96 ( .A0(n1041), .A1(n3993), .B0(n3940), .B1(n5857), .C0(n1042), 
        .Y(n667) );
  OAI221XL U97 ( .A0(n1033), .A1(n3993), .B0(n3940), .B1(n5889), .C0(n1034), 
        .Y(n665) );
  OAI221XL U98 ( .A0(n957), .A1(n3995), .B0(n3942), .B1(n5801), .C0(n958), .Y(
        n646) );
  OAI221XL U99 ( .A0(n945), .A1(n3995), .B0(n3942), .B1(n5849), .C0(n946), .Y(
        n643) );
  OAI221XL U100 ( .A0(n937), .A1(n3996), .B0(n3942), .B1(n5881), .C0(n938), 
        .Y(n641) );
  OAI221XL U101 ( .A0(n929), .A1(n3996), .B0(n3943), .B1(n5778), .C0(n930), 
        .Y(n639) );
  OAI221XL U102 ( .A0(n925), .A1(n3996), .B0(n3943), .B1(n5811), .C0(n926), 
        .Y(n638) );
  OAI221XL U103 ( .A0(n913), .A1(n3996), .B0(n3943), .B1(n5859), .C0(n914), 
        .Y(n635) );
  OAI221XL U104 ( .A0(n905), .A1(n3996), .B0(n3943), .B1(n5891), .C0(n906), 
        .Y(n633) );
  OAI221XL U105 ( .A0(n1129), .A1(n742), .B0(n3938), .B1(n5884), .C0(n1130), 
        .Y(n689) );
  OAI221XL U106 ( .A0(n1233), .A1(n3992), .B0(n3935), .B1(n5854), .C0(n1234), 
        .Y(n715) );
  OAI221XL U107 ( .A0(n1029), .A1(n3993), .B0(n3940), .B1(n5786), .C0(n1030), 
        .Y(n664) );
  OAI221XL U108 ( .A0(n1013), .A1(n3994), .B0(n3941), .B1(n5834), .C0(n1014), 
        .Y(n660) );
  OAI221XL U109 ( .A0(n885), .A1(n3997), .B0(n3944), .B1(n5832), .C0(n886), 
        .Y(n628) );
  OAI221XL U110 ( .A0(n1009), .A1(n3994), .B0(n3941), .B1(n5850), .C0(n1010), 
        .Y(n659) );
  OAI221XL U111 ( .A0(n881), .A1(n3997), .B0(n3944), .B1(n5848), .C0(n882), 
        .Y(n627) );
  OAI221XL U112 ( .A0(n1133), .A1(n742), .B0(n3938), .B1(n5868), .C0(n1134), 
        .Y(n690) );
  OAI221XL U113 ( .A0(n877), .A1(n3997), .B0(n3944), .B1(n5864), .C0(n878), 
        .Y(n626) );
  OAI221XL U114 ( .A0(n889), .A1(n3997), .B0(n3944), .B1(n5816), .C0(n890), 
        .Y(n629) );
  OAI221XL U115 ( .A0(n893), .A1(n3997), .B0(n3944), .B1(n5800), .C0(n894), 
        .Y(n630) );
  OAI221XL U116 ( .A0(n1105), .A1(n4004), .B0(n3938), .B1(n5856), .C0(n1106), 
        .Y(n683) );
  OAI221XL U117 ( .A0(n977), .A1(n3995), .B0(n3941), .B1(n5858), .C0(n978), 
        .Y(n651) );
  OAI221XL U118 ( .A0(n809), .A1(n3999), .B0(n3946), .B1(n5879), .C0(n810), 
        .Y(n609) );
  OAI221XL U119 ( .A0(n805), .A1(n3999), .B0(n3946), .B1(n5797), .C0(n806), 
        .Y(n608) );
  OAI221XL U120 ( .A0(n797), .A1(n3999), .B0(n3946), .B1(n5813), .C0(n798), 
        .Y(n606) );
  OAI221XL U121 ( .A0(n789), .A1(n3999), .B0(n3946), .B1(n5845), .C0(n790), 
        .Y(n604) );
  OAI221XL U122 ( .A0(n785), .A1(n3999), .B0(n3946), .B1(n5861), .C0(n786), 
        .Y(n603) );
  OAI221XL U123 ( .A0(n781), .A1(n3999), .B0(n3946), .B1(n5877), .C0(n782), 
        .Y(n602) );
  OAI221XL U124 ( .A0(n777), .A1(n4000), .B0(n3946), .B1(n5893), .C0(n778), 
        .Y(n601) );
  OAI221XL U125 ( .A0(n833), .A1(n3998), .B0(n3945), .B1(n5766), .C0(n834), 
        .Y(n615) );
  OAI221XL U126 ( .A0(n829), .A1(n3998), .B0(n3945), .B1(n5799), .C0(n830), 
        .Y(n614) );
  OAI221XL U127 ( .A0(n821), .A1(n3998), .B0(n3945), .B1(n5831), .C0(n822), 
        .Y(n612) );
  OAI221XL U128 ( .A0(n817), .A1(n3999), .B0(n3945), .B1(n5847), .C0(n818), 
        .Y(n611) );
  OAI221XL U129 ( .A0(n1141), .A1(n4001), .B0(n3937), .B1(n5836), .C0(n1142), 
        .Y(n692) );
  OAI221XL U130 ( .A0(n1137), .A1(n4003), .B0(n3937), .B1(n5852), .C0(n1138), 
        .Y(n691) );
  OAI221XL U131 ( .A0(n1005), .A1(n3994), .B0(n3935), .B1(n5866), .C0(n1006), 
        .Y(n658) );
  OAI221XL U132 ( .A0(n1145), .A1(n4004), .B0(n3937), .B1(n5820), .C0(n1146), 
        .Y(n693) );
  OAI221XL U133 ( .A0(n1149), .A1(n4003), .B0(n3937), .B1(n5804), .C0(n1150), 
        .Y(n694) );
  OAI221XL U134 ( .A0(n1157), .A1(n4002), .B0(n3937), .B1(n5788), .C0(n1158), 
        .Y(n696) );
  OAI221XL U135 ( .A0(n1165), .A1(n742), .B0(n3937), .B1(n5871), .C0(n1166), 
        .Y(n698) );
  OAI221XL U136 ( .A0(n1017), .A1(n3994), .B0(n3940), .B1(n5818), .C0(n1018), 
        .Y(n661) );
  OAI221XL U137 ( .A0(n1021), .A1(n3993), .B0(n3940), .B1(n5802), .C0(n1022), 
        .Y(n662) );
  OAI221XL U138 ( .A0(n901), .A1(n3996), .B0(n3943), .B1(n5784), .C0(n902), 
        .Y(n632) );
  OAI221XL U139 ( .A0(n917), .A1(n3996), .B0(n3943), .B1(n5843), .C0(n918), 
        .Y(n636) );
  OAI221XL U140 ( .A0(n1057), .A1(n3993), .B0(n3939), .B1(n5777), .C0(n1058), 
        .Y(n671) );
  OAI221XL U141 ( .A0(n753), .A1(n4000), .B0(n3947), .B1(n5846), .C0(n754), 
        .Y(n595) );
  OAI221XL U142 ( .A0(n761), .A1(n4000), .B0(n3947), .B1(n5814), .C0(n762), 
        .Y(n597) );
  OAI221XL U143 ( .A0(n765), .A1(n4000), .B0(n3947), .B1(n5798), .C0(n766), 
        .Y(n598) );
  OAI221XL U144 ( .A0(n757), .A1(n4000), .B0(n3947), .B1(n5830), .C0(n758), 
        .Y(n596) );
  OAI221XL U145 ( .A0(n749), .A1(n4000), .B0(n3947), .B1(n5862), .C0(n750), 
        .Y(n594) );
  OAI221XL U146 ( .A0(n773), .A1(n4000), .B0(n3947), .B1(n5782), .C0(n774), 
        .Y(n600) );
  OAI221XL U147 ( .A0(n1001), .A1(n3994), .B0(n3941), .B1(n5882), .C0(n1002), 
        .Y(n657) );
  OAI221XL U148 ( .A0(n873), .A1(n3997), .B0(n3944), .B1(n5880), .C0(n874), 
        .Y(n625) );
  OAI221XL U149 ( .A0(n741), .A1(n4000), .B0(n3947), .B1(n5878), .C0(n743), 
        .Y(n593) );
  OAI221XL U150 ( .A0(n1025), .A1(n3993), .B0(n3940), .B1(n5769), .C0(n1026), 
        .Y(n663) );
  XOR2X1 U151 ( .A(new_sboxw[17]), .B(n293), .Y(n5447) );
  OAI221XL U152 ( .A0(n1117), .A1(n4001), .B0(n3938), .B1(n5808), .C0(n1118), 
        .Y(n686) );
  OAI221XL U153 ( .A0(n1113), .A1(n4002), .B0(n3938), .B1(n5824), .C0(n1114), 
        .Y(n685) );
  OAI221XL U154 ( .A0(n1097), .A1(n4001), .B0(n3938), .B1(n5888), .C0(n1098), 
        .Y(n681) );
  OAI221XL U155 ( .A0(n989), .A1(n3994), .B0(n3941), .B1(n5810), .C0(n990), 
        .Y(n654) );
  OAI221XL U156 ( .A0(n985), .A1(n3994), .B0(n3941), .B1(n5826), .C0(n986), 
        .Y(n653) );
  OAI221XL U157 ( .A0(n865), .A1(n3997), .B0(n3944), .B1(n5774), .C0(n866), 
        .Y(n623) );
  OAI221XL U158 ( .A0(n861), .A1(n3997), .B0(n3944), .B1(n5812), .C0(n862), 
        .Y(n622) );
  OAI221XL U159 ( .A0(n857), .A1(n3998), .B0(n3944), .B1(n5828), .C0(n858), 
        .Y(n621) );
  OAI221XL U160 ( .A0(n801), .A1(n3999), .B0(n3946), .B1(n5776), .C0(n802), 
        .Y(n607) );
  OAI221XL U161 ( .A0(n853), .A1(n3998), .B0(n3945), .B1(n5844), .C0(n854), 
        .Y(n620) );
  OAI221XL U162 ( .A0(n849), .A1(n3998), .B0(n3945), .B1(n5860), .C0(n850), 
        .Y(n619) );
  OAI221XL U163 ( .A0(n841), .A1(n3998), .B0(n3945), .B1(n5892), .C0(n842), 
        .Y(n617) );
  OAI221XL U164 ( .A0(n1153), .A1(n4001), .B0(n3937), .B1(n5771), .C0(n1154), 
        .Y(n695) );
  OAI221XL U165 ( .A0(n1245), .A1(n3992), .B0(n3935), .B1(n5806), .C0(n1246), 
        .Y(n718) );
  OAI221XL U166 ( .A0(n1241), .A1(n3992), .B0(n3935), .B1(n5822), .C0(n1242), 
        .Y(n717) );
  OAI221XL U167 ( .A0(n1237), .A1(n3992), .B0(n3935), .B1(n5838), .C0(n1238), 
        .Y(n716) );
  OAI221XL U168 ( .A0(n1225), .A1(n3992), .B0(n3935), .B1(n5886), .C0(n1226), 
        .Y(n713) );
  OAI221XL U169 ( .A0(n897), .A1(n3997), .B0(n3943), .B1(n5770), .C0(n898), 
        .Y(n631) );
  OAI221XL U170 ( .A0(n969), .A1(n3995), .B0(n3942), .B1(n5890), .C0(n970), 
        .Y(n649) );
  OAI221XL U171 ( .A0(n1249), .A1(n3992), .B0(n3941), .B1(n5781), .C0(n1250), 
        .Y(n719) );
  OAI221XL U172 ( .A0(n1121), .A1(n4002), .B0(n3938), .B1(n5775), .C0(n1122), 
        .Y(n687) );
  OAI221XL U173 ( .A0(n1109), .A1(n4005), .B0(n3938), .B1(n5840), .C0(n1110), 
        .Y(n684) );
  OAI221XL U174 ( .A0(n993), .A1(n3994), .B0(n3941), .B1(n5780), .C0(n994), 
        .Y(n655) );
  OAI221XL U175 ( .A0(n981), .A1(n3994), .B0(n3941), .B1(n5842), .C0(n982), 
        .Y(n652) );
  OAI221XL U176 ( .A0(n769), .A1(n4000), .B0(n3947), .B1(n5768), .C0(n770), 
        .Y(n599) );
  BUFX2 U177 ( .A(n4577), .Y(n4576) );
  BUFX2 U178 ( .A(n4579), .Y(n4573) );
  BUFX2 U179 ( .A(n4579), .Y(n4572) );
  BUFX2 U180 ( .A(n4578), .Y(n4575) );
  BUFX2 U181 ( .A(n4578), .Y(n4574) );
  BUFX2 U182 ( .A(n4582), .Y(n4567) );
  BUFX2 U183 ( .A(n4582), .Y(n4566) );
  BUFX2 U184 ( .A(n4580), .Y(n4571) );
  BUFX2 U185 ( .A(n4580), .Y(n4570) );
  BUFX2 U186 ( .A(n4581), .Y(n4569) );
  BUFX2 U187 ( .A(n4581), .Y(n4568) );
  BUFX2 U188 ( .A(n4583), .Y(n4565) );
  BUFX2 U189 ( .A(n4584), .Y(n4583) );
  BUFX2 U190 ( .A(n4583), .Y(n4577) );
  BUFX2 U191 ( .A(n4585), .Y(n4579) );
  BUFX2 U192 ( .A(n4585), .Y(n4578) );
  BUFX2 U193 ( .A(n4584), .Y(n4582) );
  BUFX2 U194 ( .A(n4585), .Y(n4580) );
  BUFX2 U195 ( .A(n4584), .Y(n4581) );
  BUFX2 U196 ( .A(n4586), .Y(n4584) );
  BUFX2 U197 ( .A(n4586), .Y(n4585) );
  INVX1 U198 ( .A(reset_n), .Y(n4586) );
  INVX1 U199 ( .A(n2), .Y(n3934) );
  INVX1 U200 ( .A(n3962), .Y(n3939) );
  INVX1 U201 ( .A(n3961), .Y(n3942) );
  INVX1 U202 ( .A(n3961), .Y(n3936) );
  INVX1 U203 ( .A(n3962), .Y(n3943) );
  INVX1 U204 ( .A(n3962), .Y(n3935) );
  INVX1 U205 ( .A(n3961), .Y(n3940) );
  INVX1 U206 ( .A(n3961), .Y(n3937) );
  INVX1 U207 ( .A(n2), .Y(n3938) );
  INVX1 U208 ( .A(n3962), .Y(n3941) );
  INVX1 U209 ( .A(n3961), .Y(n3944) );
  INVX1 U210 ( .A(n3961), .Y(n3945) );
  INVX1 U211 ( .A(n3961), .Y(n3946) );
  INVX1 U212 ( .A(n3962), .Y(n3947) );
  INVX1 U213 ( .A(n3960), .Y(n1728) );
  INVX1 U214 ( .A(n3948), .Y(n1736) );
  INVX1 U215 ( .A(n3963), .Y(n3928) );
  INVX1 U216 ( .A(n3963), .Y(n3929) );
  INVX1 U217 ( .A(n3963), .Y(n3930) );
  INVX1 U218 ( .A(n3960), .Y(n3931) );
  INVX1 U219 ( .A(n3962), .Y(n3932) );
  INVX1 U220 ( .A(n3960), .Y(n3933) );
  INVX1 U221 ( .A(n3948), .Y(n1719) );
  INVX1 U222 ( .A(n3948), .Y(n1720) );
  BUFX2 U223 ( .A(n1662), .Y(n1652) );
  BUFX2 U224 ( .A(n1662), .Y(n1651) );
  BUFX2 U225 ( .A(n1661), .Y(n1653) );
  BUFX2 U226 ( .A(n1661), .Y(n1654) );
  BUFX2 U227 ( .A(n1660), .Y(n1655) );
  BUFX2 U228 ( .A(n1659), .Y(n1657) );
  BUFX2 U229 ( .A(n1660), .Y(n1656) );
  BUFX2 U230 ( .A(n1659), .Y(n1658) );
  BUFX2 U231 ( .A(n3960), .Y(n3948) );
  BUFX2 U232 ( .A(n2), .Y(n3957) );
  BUFX2 U233 ( .A(n2), .Y(n3956) );
  BUFX2 U234 ( .A(n2), .Y(n3955) );
  BUFX2 U235 ( .A(n3962), .Y(n3954) );
  BUFX2 U236 ( .A(n3962), .Y(n3953) );
  BUFX2 U237 ( .A(n3962), .Y(n3952) );
  BUFX2 U238 ( .A(n3963), .Y(n3951) );
  BUFX2 U239 ( .A(n3963), .Y(n3950) );
  BUFX2 U240 ( .A(n3963), .Y(n3949) );
  BUFX2 U241 ( .A(n5674), .Y(n1661) );
  BUFX2 U242 ( .A(n5674), .Y(n1662) );
  BUFX2 U243 ( .A(n5674), .Y(n1659) );
  BUFX2 U244 ( .A(n5674), .Y(n1660) );
  BUFX2 U245 ( .A(n1603), .Y(n1601) );
  BUFX2 U246 ( .A(n1605), .Y(n1597) );
  BUFX2 U247 ( .A(n1604), .Y(n1598) );
  BUFX2 U248 ( .A(n1604), .Y(n1599) );
  BUFX2 U249 ( .A(n1603), .Y(n1600) );
  BUFX2 U250 ( .A(n1605), .Y(n1596) );
  BUFX2 U251 ( .A(n1663), .Y(n1650) );
  BUFX2 U252 ( .A(n5674), .Y(n1663) );
  BUFX2 U253 ( .A(n2), .Y(n3962) );
  BUFX2 U254 ( .A(n2), .Y(n3963) );
  INVX1 U255 ( .A(n4220), .Y(n4203) );
  INVX1 U256 ( .A(n4253), .Y(n4231) );
  INVX1 U257 ( .A(n4219), .Y(n4204) );
  INVX1 U258 ( .A(n4254), .Y(n4232) );
  INVX1 U259 ( .A(n4218), .Y(n4205) );
  INVX1 U260 ( .A(n4252), .Y(n4233) );
  INVX1 U261 ( .A(n4217), .Y(n4206) );
  INVX1 U262 ( .A(n4251), .Y(n4234) );
  INVX1 U263 ( .A(n4252), .Y(n4235) );
  INVX1 U264 ( .A(n4215), .Y(n4207) );
  INVX1 U265 ( .A(n4251), .Y(n4236) );
  INVX1 U266 ( .A(n4220), .Y(n4208) );
  INVX1 U267 ( .A(n4250), .Y(n4237) );
  INVX1 U268 ( .A(n4219), .Y(n4209) );
  INVX1 U269 ( .A(n4249), .Y(n4238) );
  INVX1 U270 ( .A(n4217), .Y(n4210) );
  INVX1 U271 ( .A(n4248), .Y(n4239) );
  INVX1 U272 ( .A(n4218), .Y(n4211) );
  INVX1 U273 ( .A(n4247), .Y(n4240) );
  INVX1 U274 ( .A(n4215), .Y(n4212) );
  INVX1 U275 ( .A(n4246), .Y(n4241) );
  INVX1 U276 ( .A(n4214), .Y(n4213) );
  INVX1 U277 ( .A(n4245), .Y(n4242) );
  BUFX2 U278 ( .A(n1617), .Y(n1615) );
  BUFX2 U279 ( .A(n1618), .Y(n1614) );
  BUFX2 U280 ( .A(n1620), .Y(n1610) );
  BUFX2 U281 ( .A(n1619), .Y(n1611) );
  BUFX2 U282 ( .A(n1619), .Y(n1612) );
  BUFX2 U283 ( .A(n1618), .Y(n1613) );
  BUFX2 U284 ( .A(n1617), .Y(n1616) );
  BUFX2 U285 ( .A(n1620), .Y(n1609) );
  BUFX2 U286 ( .A(n5668), .Y(n1602) );
  BUFX2 U287 ( .A(n5668), .Y(n1606) );
  BUFX2 U288 ( .A(n5668), .Y(n1605) );
  BUFX2 U289 ( .A(n5668), .Y(n1604) );
  BUFX2 U290 ( .A(n5668), .Y(n1603) );
  BUFX2 U291 ( .A(n1645), .Y(n1643) );
  BUFX2 U292 ( .A(n1645), .Y(n1642) );
  BUFX2 U293 ( .A(n1645), .Y(n1641) );
  BUFX2 U294 ( .A(n1579), .Y(n1571) );
  BUFX2 U295 ( .A(n1646), .Y(n1640) );
  BUFX2 U296 ( .A(n1646), .Y(n1639) );
  BUFX2 U297 ( .A(n1647), .Y(n1638) );
  BUFX2 U298 ( .A(n1647), .Y(n1637) );
  BUFX2 U299 ( .A(n1607), .Y(n1595) );
  BUFX2 U300 ( .A(n5668), .Y(n1607) );
  BUFX2 U301 ( .A(n1579), .Y(n1572) );
  BUFX2 U302 ( .A(n1673), .Y(n1672) );
  BUFX2 U303 ( .A(n1676), .Y(n1667) );
  BUFX2 U304 ( .A(n1676), .Y(n1668) );
  BUFX2 U305 ( .A(n1674), .Y(n1669) );
  BUFX2 U306 ( .A(n1674), .Y(n1670) );
  BUFX2 U307 ( .A(n1673), .Y(n1671) );
  BUFX2 U308 ( .A(n1578), .Y(n1574) );
  BUFX2 U309 ( .A(n1578), .Y(n1573) );
  BUFX2 U310 ( .A(n1577), .Y(n1576) );
  BUFX2 U311 ( .A(n1577), .Y(n1575) );
  BUFX2 U312 ( .A(n1362), .Y(n1416) );
  BUFX2 U313 ( .A(n1356), .Y(n1408) );
  BUFX2 U314 ( .A(n1362), .Y(n1391) );
  BUFX2 U315 ( .A(n1358), .Y(n1401) );
  BUFX2 U316 ( .A(n1356), .Y(n1409) );
  BUFX2 U317 ( .A(n1357), .Y(n1406) );
  BUFX2 U318 ( .A(n1361), .Y(n1392) );
  BUFX2 U319 ( .A(n1356), .Y(n1407) );
  BUFX2 U320 ( .A(n1361), .Y(n1393) );
  BUFX2 U321 ( .A(n1357), .Y(n1405) );
  BUFX2 U322 ( .A(n1357), .Y(n1404) );
  BUFX2 U323 ( .A(n1354), .Y(n1413) );
  BUFX2 U324 ( .A(n1361), .Y(n1394) );
  BUFX2 U325 ( .A(n1358), .Y(n1403) );
  BUFX2 U326 ( .A(n1354), .Y(n1414) );
  BUFX2 U327 ( .A(n1360), .Y(n1395) );
  BUFX2 U328 ( .A(n1355), .Y(n1411) );
  BUFX2 U329 ( .A(n1354), .Y(n1415) );
  BUFX2 U330 ( .A(n1365), .Y(n1381) );
  BUFX2 U331 ( .A(n1355), .Y(n1410) );
  BUFX2 U332 ( .A(n1363), .Y(n1388) );
  BUFX2 U333 ( .A(n1362), .Y(n1389) );
  BUFX2 U334 ( .A(n1362), .Y(n1390) );
  BUFX2 U335 ( .A(n1358), .Y(n1402) );
  BUFX2 U336 ( .A(n1359), .Y(n1399) );
  BUFX2 U337 ( .A(n1359), .Y(n1400) );
  BUFX2 U338 ( .A(n1363), .Y(n1386) );
  BUFX2 U339 ( .A(n1365), .Y(n1382) );
  BUFX2 U340 ( .A(n1364), .Y(n1383) );
  BUFX2 U341 ( .A(n1364), .Y(n1385) );
  BUFX2 U342 ( .A(n1364), .Y(n1384) );
  BUFX2 U343 ( .A(n1360), .Y(n1396) );
  BUFX2 U344 ( .A(n1363), .Y(n1387) );
  BUFX2 U345 ( .A(n1359), .Y(n1398) );
  BUFX2 U346 ( .A(n1360), .Y(n1397) );
  BUFX2 U347 ( .A(n1355), .Y(n1412) );
  BUFX2 U348 ( .A(n1365), .Y(n1380) );
  BUFX2 U349 ( .A(n1367), .Y(n1375) );
  BUFX2 U350 ( .A(n1367), .Y(n1376) );
  BUFX2 U351 ( .A(n1366), .Y(n1378) );
  BUFX2 U352 ( .A(n1368), .Y(n1371) );
  BUFX2 U353 ( .A(n1368), .Y(n1372) );
  BUFX2 U354 ( .A(n1367), .Y(n1374) );
  BUFX2 U355 ( .A(n1366), .Y(n1377) );
  BUFX2 U356 ( .A(n1368), .Y(n1373) );
  BUFX2 U357 ( .A(n1366), .Y(n1379) );
  BUFX2 U358 ( .A(n1300), .Y(n1338) );
  BUFX2 U359 ( .A(n1300), .Y(n1337) );
  BUFX2 U360 ( .A(n1299), .Y(n1340) );
  BUFX2 U361 ( .A(n1299), .Y(n1342) );
  BUFX2 U362 ( .A(n1300), .Y(n1339) );
  BUFX2 U363 ( .A(n1301), .Y(n1335) );
  BUFX2 U364 ( .A(n1298), .Y(n1345) );
  BUFX2 U365 ( .A(n1298), .Y(n1343) );
  BUFX2 U366 ( .A(n1298), .Y(n1344) );
  BUFX2 U367 ( .A(n1301), .Y(n1336) );
  BUFX2 U368 ( .A(n1301), .Y(n1334) );
  BUFX2 U369 ( .A(n1299), .Y(n1341) );
  BUFX2 U370 ( .A(n1304), .Y(n1328) );
  BUFX2 U371 ( .A(n1306), .Y(n1317) );
  BUFX2 U372 ( .A(n1304), .Y(n1321) );
  BUFX2 U373 ( .A(n1307), .Y(n1322) );
  BUFX2 U374 ( .A(n1294), .Y(n1323) );
  BUFX2 U375 ( .A(n1306), .Y(n1316) );
  BUFX2 U376 ( .A(n1307), .Y(n1313) );
  BUFX2 U377 ( .A(n1307), .Y(n1312) );
  BUFX2 U378 ( .A(n1302), .Y(n1331) );
  BUFX2 U379 ( .A(n1300), .Y(n1329) );
  BUFX2 U380 ( .A(n1296), .Y(n1330) );
  BUFX2 U381 ( .A(n1302), .Y(n1333) );
  BUFX2 U382 ( .A(n1302), .Y(n1332) );
  BUFX2 U383 ( .A(n1304), .Y(n1326) );
  BUFX2 U384 ( .A(n1304), .Y(n1325) );
  BUFX2 U385 ( .A(n1304), .Y(n1324) );
  BUFX2 U386 ( .A(n1307), .Y(n1314) );
  BUFX2 U387 ( .A(n1305), .Y(n1320) );
  BUFX2 U388 ( .A(n1305), .Y(n1319) );
  BUFX2 U389 ( .A(n1305), .Y(n1318) );
  BUFX2 U390 ( .A(n1303), .Y(n1327) );
  BUFX2 U391 ( .A(n1306), .Y(n1315) );
  BUFX2 U392 ( .A(n1308), .Y(n1311) );
  BUFX2 U393 ( .A(n1308), .Y(n1310) );
  BUFX2 U394 ( .A(n1700), .Y(n1697) );
  BUFX2 U395 ( .A(n1701), .Y(n1695) );
  BUFX2 U396 ( .A(n1703), .Y(n1694) );
  BUFX2 U397 ( .A(n1702), .Y(n1693) );
  BUFX2 U398 ( .A(n1702), .Y(n1692) );
  BUFX2 U399 ( .A(n1701), .Y(n1696) );
  BUFX2 U400 ( .A(n1700), .Y(n1698) );
  BUFX2 U401 ( .A(n1308), .Y(n1309) );
  BUFX2 U402 ( .A(n4227), .Y(n4220) );
  BUFX2 U403 ( .A(n4254), .Y(n4253) );
  BUFX2 U404 ( .A(n4227), .Y(n4219) );
  BUFX2 U405 ( .A(n4227), .Y(n4218) );
  BUFX2 U406 ( .A(n4228), .Y(n4217) );
  BUFX2 U407 ( .A(n4228), .Y(n4216) );
  BUFX2 U408 ( .A(n730), .Y(n4252) );
  BUFX2 U409 ( .A(n4228), .Y(n4215) );
  BUFX2 U410 ( .A(n4230), .Y(n4251) );
  BUFX2 U411 ( .A(n4255), .Y(n4250) );
  BUFX2 U412 ( .A(n4255), .Y(n4249) );
  BUFX2 U413 ( .A(n4255), .Y(n4248) );
  BUFX2 U414 ( .A(n4256), .Y(n4247) );
  BUFX2 U415 ( .A(n4256), .Y(n4246) );
  BUFX2 U416 ( .A(n4227), .Y(n4214) );
  BUFX2 U417 ( .A(n4256), .Y(n4245) );
  BUFX2 U418 ( .A(n3961), .Y(n3959) );
  BUFX2 U419 ( .A(n3961), .Y(n3958) );
  BUFX2 U420 ( .A(n4226), .Y(n4221) );
  BUFX2 U421 ( .A(n4226), .Y(n4222) );
  BUFX2 U422 ( .A(n4226), .Y(n4223) );
  INVX1 U423 ( .A(n4333), .Y(n4314) );
  INVX1 U424 ( .A(n4365), .Y(n4342) );
  INVX1 U425 ( .A(n4332), .Y(n4315) );
  INVX1 U426 ( .A(n4365), .Y(n4343) );
  INVX1 U427 ( .A(n4335), .Y(n4316) );
  INVX1 U428 ( .A(n4364), .Y(n4344) );
  INVX1 U429 ( .A(n4335), .Y(n4317) );
  INVX1 U430 ( .A(n4363), .Y(n4345) );
  INVX1 U431 ( .A(n4334), .Y(n4318) );
  INVX1 U432 ( .A(n4362), .Y(n4346) );
  INVX1 U433 ( .A(n4333), .Y(n4319) );
  INVX1 U434 ( .A(n4361), .Y(n4347) );
  INVX1 U435 ( .A(n4332), .Y(n4320) );
  INVX1 U436 ( .A(n4360), .Y(n4348) );
  INVX1 U437 ( .A(n4331), .Y(n4321) );
  INVX1 U438 ( .A(n4359), .Y(n4349) );
  INVX1 U439 ( .A(n4330), .Y(n4322) );
  INVX1 U440 ( .A(n4358), .Y(n4350) );
  INVX1 U441 ( .A(n4329), .Y(n4323) );
  INVX1 U442 ( .A(n4357), .Y(n4351) );
  INVX1 U443 ( .A(n4328), .Y(n4324) );
  INVX1 U444 ( .A(n4356), .Y(n4352) );
  INVX1 U445 ( .A(n4327), .Y(n4325) );
  INVX1 U446 ( .A(n4355), .Y(n4353) );
  BUFX2 U447 ( .A(n4227), .Y(n4224) );
  BUFX2 U448 ( .A(n4229), .Y(n4225) );
  INVX1 U449 ( .A(n4244), .Y(n4243) );
  BUFX2 U450 ( .A(n3961), .Y(n3960) );
  INVXL U451 ( .A(new_sboxw[11]), .Y(n5220) );
  INVXL U452 ( .A(new_sboxw[15]), .Y(n5351) );
  INVXL U453 ( .A(new_sboxw[1]), .Y(n4891) );
  BUFX2 U454 ( .A(n5669), .Y(n1617) );
  BUFX2 U455 ( .A(n5669), .Y(n1620) );
  BUFX2 U456 ( .A(n5669), .Y(n1619) );
  BUFX2 U457 ( .A(n5669), .Y(n1618) );
  BUFX2 U458 ( .A(n1621), .Y(n1608) );
  BUFX2 U459 ( .A(n5669), .Y(n1621) );
  NAND2BX1 U460 ( .AN(n3992), .B(n4544), .Y(n4603) );
  BUFX2 U461 ( .A(n5672), .Y(n1648) );
  BUFX2 U462 ( .A(n5672), .Y(n1644) );
  BUFX2 U463 ( .A(n5672), .Y(n1645) );
  BUFX2 U464 ( .A(n5672), .Y(n1646) );
  BUFX2 U465 ( .A(n5672), .Y(n1647) );
  BUFX2 U466 ( .A(n1568), .Y(n1578) );
  BUFX2 U467 ( .A(n1664), .Y(n1676) );
  BUFX2 U468 ( .A(n1665), .Y(n1675) );
  BUFX2 U469 ( .A(n1664), .Y(n1674) );
  BUFX2 U470 ( .A(n1568), .Y(n1577) );
  BUFX2 U471 ( .A(n1664), .Y(n1673) );
  BUFX2 U472 ( .A(n1568), .Y(n1579) );
  BUFX2 U473 ( .A(n1634), .Y(n1623) );
  BUFX2 U474 ( .A(n1633), .Y(n1625) );
  BUFX2 U475 ( .A(n1563), .Y(n1558) );
  BUFX2 U476 ( .A(n1649), .Y(n1636) );
  BUFX2 U477 ( .A(n5672), .Y(n1649) );
  BUFX2 U478 ( .A(n1563), .Y(n1559) );
  BUFX2 U479 ( .A(n1631), .Y(n1630) );
  BUFX2 U480 ( .A(n1635), .Y(n1624) );
  BUFX2 U481 ( .A(n1633), .Y(n1626) );
  BUFX2 U482 ( .A(n1632), .Y(n1627) );
  BUFX2 U483 ( .A(n1632), .Y(n1628) );
  BUFX2 U484 ( .A(n1631), .Y(n1629) );
  BUFX2 U485 ( .A(n1562), .Y(n1560) );
  BUFX2 U486 ( .A(n1590), .Y(n1588) );
  BUFX2 U487 ( .A(n1591), .Y(n1587) );
  BUFX2 U488 ( .A(n1594), .Y(n1582) );
  BUFX2 U489 ( .A(n1593), .Y(n1583) );
  BUFX2 U490 ( .A(n1592), .Y(n1584) );
  BUFX2 U491 ( .A(n1592), .Y(n1585) );
  BUFX2 U492 ( .A(n1591), .Y(n1586) );
  BUFX2 U493 ( .A(n1562), .Y(n1561) );
  BUFX2 U494 ( .A(n1590), .Y(n1589) );
  BUFX2 U495 ( .A(n1266), .Y(n1275) );
  BUFX2 U496 ( .A(n1268), .Y(n1271) );
  BUFX2 U497 ( .A(n1266), .Y(n1274) );
  BUFX2 U498 ( .A(n1351), .Y(n1362) );
  BUFX2 U499 ( .A(n1353), .Y(n1356) );
  BUFX2 U500 ( .A(n1295), .Y(n1300) );
  BUFX2 U501 ( .A(n1352), .Y(n1357) );
  BUFX2 U502 ( .A(n1351), .Y(n1361) );
  BUFX2 U503 ( .A(n1293), .Y(n1306) );
  BUFX2 U504 ( .A(n1352), .Y(n1358) );
  BUFX2 U505 ( .A(n1353), .Y(n1354) );
  BUFX2 U506 ( .A(n1296), .Y(n1299) );
  BUFX2 U507 ( .A(n1353), .Y(n1355) );
  BUFX2 U508 ( .A(n1295), .Y(n1302) );
  BUFX2 U509 ( .A(n1294), .Y(n1304) );
  BUFX2 U510 ( .A(n1293), .Y(n1307) );
  BUFX2 U511 ( .A(n1350), .Y(n1365) );
  BUFX2 U512 ( .A(n1296), .Y(n1298) );
  BUFX2 U513 ( .A(n1350), .Y(n1364) );
  BUFX2 U514 ( .A(n1294), .Y(n1305) );
  BUFX2 U515 ( .A(n1349), .Y(n1367) );
  BUFX2 U516 ( .A(n1349), .Y(n1366) );
  BUFX2 U517 ( .A(n1295), .Y(n1301) );
  BUFX2 U518 ( .A(n1350), .Y(n1363) );
  BUFX2 U519 ( .A(n1352), .Y(n1359) );
  BUFX2 U520 ( .A(n1349), .Y(n1368) );
  BUFX2 U521 ( .A(n1351), .Y(n1360) );
  BUFX2 U522 ( .A(n1293), .Y(n1303) );
  BUFX2 U523 ( .A(n1293), .Y(n1308) );
  BUFX2 U524 ( .A(n1353), .Y(n1369) );
  BUFX2 U525 ( .A(n1418), .Y(n1370) );
  BUFX2 U526 ( .A(n1297), .Y(n1346) );
  BUFX2 U527 ( .A(n1296), .Y(n1297) );
  BUFX2 U528 ( .A(n1565), .Y(n1554) );
  BUFX2 U529 ( .A(n1565), .Y(n1555) );
  BUFX2 U530 ( .A(n1565), .Y(n1557) );
  BUFX2 U531 ( .A(n1564), .Y(n1556) );
  BUFX2 U532 ( .A(n1268), .Y(n1270) );
  BUFX2 U533 ( .A(n1267), .Y(n1272) );
  BUFX2 U534 ( .A(n1267), .Y(n1273) );
  BUFX2 U535 ( .A(n1688), .Y(n1682) );
  BUFX2 U536 ( .A(n1687), .Y(n1683) );
  BUFX2 U537 ( .A(n5758), .Y(n1699) );
  BUFX2 U538 ( .A(n5758), .Y(n1702) );
  BUFX2 U539 ( .A(n1281), .Y(n1285) );
  BUFX2 U540 ( .A(n1282), .Y(n1284) );
  BUFX2 U541 ( .A(n1280), .Y(n1287) );
  BUFX2 U542 ( .A(n1280), .Y(n1288) );
  BUFX2 U543 ( .A(n1281), .Y(n1286) );
  BUFX2 U544 ( .A(n5758), .Y(n1700) );
  BUFX2 U545 ( .A(n5758), .Y(n1701) );
  BUFX2 U546 ( .A(n1282), .Y(n1283) );
  BUFX2 U547 ( .A(n1703), .Y(n1691) );
  BUFX2 U548 ( .A(n5758), .Y(n1703) );
  BUFX2 U549 ( .A(n1689), .Y(n1680) );
  BUFX2 U550 ( .A(n1689), .Y(n1679) );
  BUFX2 U551 ( .A(n1688), .Y(n1681) );
  BUFX2 U552 ( .A(n1687), .Y(n1684) );
  BUFX2 U553 ( .A(n1713), .Y(n1710) );
  BUFX2 U554 ( .A(n1714), .Y(n1708) );
  BUFX2 U555 ( .A(n4003), .Y(n3995) );
  BUFX2 U556 ( .A(n4004), .Y(n3993) );
  BUFX2 U557 ( .A(n4003), .Y(n3996) );
  BUFX2 U558 ( .A(n1715), .Y(n1707) );
  BUFX2 U559 ( .A(n1715), .Y(n1706) );
  BUFX2 U560 ( .A(n1716), .Y(n1705) );
  BUFX2 U561 ( .A(n1716), .Y(n1704) );
  BUFX2 U562 ( .A(n1714), .Y(n1709) );
  BUFX2 U563 ( .A(n1715), .Y(n1712) );
  BUFX2 U564 ( .A(n1713), .Y(n1711) );
  BUFX2 U565 ( .A(n4004), .Y(n3994) );
  BUFX2 U566 ( .A(n4002), .Y(n3997) );
  BUFX2 U567 ( .A(n4002), .Y(n3998) );
  BUFX2 U568 ( .A(n4001), .Y(n3999) );
  BUFX2 U569 ( .A(n4001), .Y(n4000) );
  BUFX2 U570 ( .A(n4257), .Y(n4244) );
  BUFX2 U571 ( .A(n4230), .Y(n4257) );
  BUFX2 U572 ( .A(n722), .Y(n4365) );
  BUFX2 U573 ( .A(n722), .Y(n4364) );
  BUFX2 U574 ( .A(n4339), .Y(n4335) );
  BUFX2 U575 ( .A(n4367), .Y(n4363) );
  BUFX2 U576 ( .A(n4339), .Y(n4334) );
  BUFX2 U577 ( .A(n4367), .Y(n4362) );
  BUFX2 U578 ( .A(n4339), .Y(n4333) );
  BUFX2 U579 ( .A(n4367), .Y(n4361) );
  BUFX2 U580 ( .A(n4340), .Y(n4332) );
  BUFX2 U581 ( .A(n4368), .Y(n4360) );
  BUFX2 U582 ( .A(n4368), .Y(n4359) );
  BUFX2 U583 ( .A(n4340), .Y(n4330) );
  BUFX2 U584 ( .A(n4368), .Y(n4358) );
  BUFX2 U585 ( .A(n4341), .Y(n4329) );
  BUFX2 U586 ( .A(n4369), .Y(n4357) );
  BUFX2 U587 ( .A(n4369), .Y(n4356) );
  BUFX2 U588 ( .A(n4341), .Y(n4327) );
  BUFX2 U589 ( .A(n4340), .Y(n4331) );
  BUFX2 U590 ( .A(n4341), .Y(n4328) );
  BUFX2 U591 ( .A(n4369), .Y(n4355) );
  BUFX2 U592 ( .A(n4229), .Y(n4226) );
  BUFX2 U593 ( .A(n4338), .Y(n4337) );
  BUFX2 U594 ( .A(n2), .Y(n3961) );
  BUFX2 U595 ( .A(n5761), .Y(n1717) );
  BUFX2 U596 ( .A(n722), .Y(n4366) );
  INVX1 U597 ( .A(n4110), .Y(n4094) );
  INVX1 U598 ( .A(n3988), .Y(n3964) );
  INVX1 U599 ( .A(n3987), .Y(n3965) );
  INVX1 U600 ( .A(n3986), .Y(n3966) );
  INVX1 U601 ( .A(n3985), .Y(n3967) );
  INVX1 U602 ( .A(n3984), .Y(n3968) );
  INVX1 U603 ( .A(n3983), .Y(n3969) );
  INVX1 U604 ( .A(n3982), .Y(n3970) );
  INVX1 U605 ( .A(n3981), .Y(n3971) );
  INVX1 U606 ( .A(n3980), .Y(n3972) );
  INVX1 U607 ( .A(n3979), .Y(n3973) );
  INVX1 U608 ( .A(n3978), .Y(n3974) );
  INVX1 U609 ( .A(n3977), .Y(n3975) );
  INVX1 U610 ( .A(n4029), .Y(n4006) );
  INVX1 U611 ( .A(n4053), .Y(n4034) );
  INVX1 U612 ( .A(n4086), .Y(n4062) );
  INVX1 U613 ( .A(n4114), .Y(n4090) );
  INVX1 U614 ( .A(n4142), .Y(n4118) );
  INVX1 U615 ( .A(n4170), .Y(n4146) );
  INVX1 U616 ( .A(n4198), .Y(n4174) );
  INVX1 U617 ( .A(n4282), .Y(n4258) );
  INVX1 U618 ( .A(n727), .Y(n4286) );
  INVX1 U619 ( .A(n4028), .Y(n4007) );
  INVX1 U620 ( .A(n4055), .Y(n4035) );
  INVX1 U621 ( .A(n4086), .Y(n4063) );
  INVX1 U622 ( .A(n4113), .Y(n4091) );
  INVX1 U623 ( .A(n4141), .Y(n4119) );
  INVX1 U624 ( .A(n4169), .Y(n4147) );
  INVX1 U625 ( .A(n4197), .Y(n4175) );
  INVX1 U626 ( .A(n4281), .Y(n4259) );
  INVX1 U627 ( .A(n4309), .Y(n4287) );
  INVX1 U628 ( .A(n4027), .Y(n4008) );
  INVX1 U629 ( .A(n4056), .Y(n4036) );
  INVX1 U630 ( .A(n4077), .Y(n4064) );
  INVX1 U631 ( .A(n4112), .Y(n4092) );
  INVX1 U632 ( .A(n4140), .Y(n4120) );
  INVX1 U633 ( .A(n4168), .Y(n4148) );
  INVX1 U634 ( .A(n4196), .Y(n4176) );
  INVX1 U635 ( .A(n4280), .Y(n4260) );
  INVX1 U636 ( .A(n4308), .Y(n4288) );
  INVX1 U637 ( .A(n4026), .Y(n4009) );
  INVX1 U638 ( .A(n4055), .Y(n4037) );
  INVX1 U639 ( .A(n4083), .Y(n4065) );
  INVX1 U640 ( .A(n4111), .Y(n4093) );
  INVX1 U641 ( .A(n4139), .Y(n4121) );
  INVX1 U642 ( .A(n4167), .Y(n4149) );
  INVX1 U643 ( .A(n4195), .Y(n4177) );
  INVX1 U644 ( .A(n4279), .Y(n4261) );
  INVX1 U645 ( .A(n4307), .Y(n4289) );
  INVX1 U646 ( .A(n4026), .Y(n4010) );
  INVX1 U647 ( .A(n4054), .Y(n4038) );
  INVX1 U648 ( .A(n4082), .Y(n4066) );
  INVX1 U649 ( .A(n4138), .Y(n4122) );
  INVX1 U650 ( .A(n4166), .Y(n4150) );
  INVX1 U651 ( .A(n4194), .Y(n4178) );
  INVX1 U652 ( .A(n4278), .Y(n4262) );
  INVX1 U653 ( .A(n4306), .Y(n4290) );
  INVX1 U654 ( .A(n4025), .Y(n4011) );
  INVX1 U655 ( .A(n4053), .Y(n4039) );
  INVX1 U656 ( .A(n4081), .Y(n4067) );
  INVX1 U657 ( .A(n4109), .Y(n4095) );
  INVX1 U658 ( .A(n4137), .Y(n4123) );
  INVX1 U659 ( .A(n4165), .Y(n4151) );
  INVX1 U660 ( .A(n4193), .Y(n4179) );
  INVX1 U661 ( .A(n4277), .Y(n4263) );
  INVX1 U662 ( .A(n4305), .Y(n4291) );
  INVX1 U663 ( .A(n4024), .Y(n4012) );
  INVX1 U664 ( .A(n4052), .Y(n4040) );
  INVX1 U665 ( .A(n4080), .Y(n4068) );
  INVX1 U666 ( .A(n4108), .Y(n4096) );
  INVX1 U667 ( .A(n4136), .Y(n4124) );
  INVX1 U668 ( .A(n4164), .Y(n4152) );
  INVX1 U669 ( .A(n4192), .Y(n4180) );
  INVX1 U670 ( .A(n4276), .Y(n4264) );
  INVX1 U671 ( .A(n4304), .Y(n4292) );
  INVX1 U672 ( .A(n4023), .Y(n4013) );
  INVX1 U673 ( .A(n4051), .Y(n4041) );
  INVX1 U674 ( .A(n4079), .Y(n4069) );
  INVX1 U675 ( .A(n4107), .Y(n4097) );
  INVX1 U676 ( .A(n4135), .Y(n4125) );
  INVX1 U677 ( .A(n4163), .Y(n4153) );
  INVX1 U678 ( .A(n4191), .Y(n4181) );
  INVX1 U679 ( .A(n4275), .Y(n4265) );
  INVX1 U680 ( .A(n4303), .Y(n4293) );
  INVX1 U681 ( .A(n4022), .Y(n4014) );
  INVX1 U682 ( .A(n4050), .Y(n4042) );
  INVX1 U683 ( .A(n4078), .Y(n4070) );
  INVX1 U684 ( .A(n4106), .Y(n4098) );
  INVX1 U685 ( .A(n4134), .Y(n4126) );
  INVX1 U686 ( .A(n4162), .Y(n4154) );
  INVX1 U687 ( .A(n4190), .Y(n4182) );
  INVX1 U688 ( .A(n4274), .Y(n4266) );
  INVX1 U689 ( .A(n4302), .Y(n4294) );
  INVX1 U690 ( .A(n4021), .Y(n4015) );
  INVX1 U691 ( .A(n4049), .Y(n4043) );
  INVX1 U692 ( .A(n4077), .Y(n4071) );
  INVX1 U693 ( .A(n4105), .Y(n4099) );
  INVX1 U694 ( .A(n4133), .Y(n4127) );
  INVX1 U695 ( .A(n4161), .Y(n4155) );
  INVX1 U696 ( .A(n4189), .Y(n4183) );
  INVX1 U697 ( .A(n4273), .Y(n4267) );
  INVX1 U698 ( .A(n4301), .Y(n4295) );
  INVX1 U699 ( .A(n4020), .Y(n4016) );
  INVX1 U700 ( .A(n4048), .Y(n4044) );
  INVX1 U701 ( .A(n4076), .Y(n4072) );
  INVX1 U702 ( .A(n4104), .Y(n4100) );
  INVX1 U703 ( .A(n4132), .Y(n4128) );
  INVX1 U704 ( .A(n4160), .Y(n4156) );
  INVX1 U705 ( .A(n4188), .Y(n4184) );
  INVX1 U706 ( .A(n4272), .Y(n4268) );
  INVX1 U707 ( .A(n4300), .Y(n4296) );
  INVX1 U708 ( .A(n4019), .Y(n4017) );
  INVX1 U709 ( .A(n4047), .Y(n4045) );
  INVX1 U710 ( .A(n4075), .Y(n4073) );
  INVX1 U711 ( .A(n4103), .Y(n4101) );
  INVX1 U712 ( .A(n4131), .Y(n4129) );
  INVX1 U713 ( .A(n4159), .Y(n4157) );
  INVX1 U714 ( .A(n4187), .Y(n4185) );
  INVX1 U715 ( .A(n4271), .Y(n4269) );
  INVX1 U716 ( .A(n4299), .Y(n4297) );
  BUFX2 U717 ( .A(n4338), .Y(n4336) );
  BUFX2 U718 ( .A(n4230), .Y(n4254) );
  BUFX2 U719 ( .A(n4229), .Y(n4227) );
  BUFX2 U720 ( .A(n4229), .Y(n4228) );
  BUFX2 U721 ( .A(n4230), .Y(n4255) );
  BUFX2 U722 ( .A(n4230), .Y(n4256) );
  INVX1 U723 ( .A(n4338), .Y(n4326) );
  INVX1 U724 ( .A(n4361), .Y(n4354) );
  INVX1 U725 ( .A(n825), .Y(n4958) );
  INVXL U726 ( .A(new_sboxw[6]), .Y(n5056) );
  INVXL U727 ( .A(new_sboxw[0]), .Y(n4858) );
  INVX1 U728 ( .A(n869), .Y(n4604) );
  BUFX2 U729 ( .A(n642), .Y(n1503) );
  INVXL U730 ( .A(new_sboxw[7]), .Y(n5088) );
  INVXL U731 ( .A(new_sboxw[13]), .Y(n5286) );
  INVXL U732 ( .A(new_sboxw[8]), .Y(n5121) );
  INVXL U733 ( .A(new_sboxw[12]), .Y(n5253) );
  INVXL U734 ( .A(new_sboxw[4]), .Y(n4990) );
  INVXL U735 ( .A(new_sboxw[2]), .Y(n4924) );
  INVXL U736 ( .A(new_sboxw[3]), .Y(n4957) );
  INVXL U737 ( .A(new_sboxw[5]), .Y(n5023) );
  INVXL U738 ( .A(new_sboxw[10]), .Y(n5187) );
  INVXL U739 ( .A(new_sboxw[14]), .Y(n5319) );
  INVX1 U740 ( .A(new_sboxw[28]), .Y(n5527) );
  INVX1 U741 ( .A(new_sboxw[30]), .Y(n5599) );
  INVX1 U742 ( .A(new_sboxw[24]), .Y(n5383) );
  INVX1 U743 ( .A(new_sboxw[25]), .Y(n5419) );
  INVX1 U744 ( .A(new_sboxw[26]), .Y(n5455) );
  INVX1 U745 ( .A(new_sboxw[27]), .Y(n5491) );
  INVX1 U746 ( .A(new_sboxw[29]), .Y(n5563) );
  INVX1 U747 ( .A(new_sboxw[31]), .Y(n5635) );
  BUFX2 U748 ( .A(n666), .Y(n1479) );
  INVX1 U749 ( .A(n861), .Y(n4667) );
  INVX1 U750 ( .A(n857), .Y(n4699) );
  INVX1 U751 ( .A(n849), .Y(n4763) );
  INVX1 U752 ( .A(n841), .Y(n4826) );
  INVX1 U753 ( .A(n829), .Y(n4925) );
  INVX1 U754 ( .A(n817), .Y(n5024) );
  INVX1 U755 ( .A(n809), .Y(n5089) );
  INVX1 U756 ( .A(n833), .Y(n4892) );
  INVX1 U757 ( .A(n5448), .Y(n899) );
  INVX1 U758 ( .A(n5556), .Y(n887) );
  INVX1 U759 ( .A(n5592), .Y(n883) );
  INVX1 U760 ( .A(n5628), .Y(n879) );
  INVX1 U761 ( .A(n5520), .Y(n891) );
  INVX1 U762 ( .A(n5484), .Y(n895) );
  INVX1 U763 ( .A(n5412), .Y(n903) );
  INVX1 U764 ( .A(n777), .Y(n5352) );
  NAND3BX1 U765 ( .AN(n4602), .B(n1714), .C(n4417), .Y(n4599) );
  INVX1 U766 ( .A(n1141), .Y(n5558) );
  INVX1 U767 ( .A(n1013), .Y(n5545) );
  INVX1 U768 ( .A(n885), .Y(n5535) );
  INVX1 U769 ( .A(n1153), .Y(n5450) );
  INVX1 U770 ( .A(n1025), .Y(n5437) );
  INVX1 U771 ( .A(n897), .Y(n5427) );
  INVX1 U772 ( .A(n1133), .Y(n5630) );
  INVX1 U773 ( .A(n1005), .Y(n5617) );
  INVX1 U774 ( .A(n877), .Y(n5607) );
  INVX1 U775 ( .A(n1157), .Y(n5414) );
  INVX1 U776 ( .A(n1029), .Y(n5401) );
  INVX1 U777 ( .A(n901), .Y(n5391) );
  INVX1 U778 ( .A(n789), .Y(n5254) );
  INVX1 U779 ( .A(n781), .Y(n5320) );
  INVX1 U780 ( .A(n805), .Y(n5122) );
  INVX1 U781 ( .A(n801), .Y(n5155) );
  INVX1 U782 ( .A(n1137), .Y(n5594) );
  INVX1 U783 ( .A(n1009), .Y(n5581) );
  INVX1 U784 ( .A(n881), .Y(n5571) );
  INVX1 U785 ( .A(n1145), .Y(n5522) );
  INVX1 U786 ( .A(n1017), .Y(n5509) );
  INVX1 U787 ( .A(n889), .Y(n5499) );
  INVX1 U788 ( .A(n1149), .Y(n5486) );
  INVX1 U789 ( .A(n1021), .Y(n5473) );
  INVX1 U790 ( .A(n893), .Y(n5463) );
  BUFX2 U791 ( .A(n5663), .Y(n1590) );
  BUFX2 U792 ( .A(n5663), .Y(n1593) );
  BUFX2 U793 ( .A(n5663), .Y(n1592) );
  BUFX2 U794 ( .A(n5663), .Y(n1591) );
  INVX1 U795 ( .A(n797), .Y(n5188) );
  INVX1 U796 ( .A(n793), .Y(n5221) );
  INVX1 U797 ( .A(n785), .Y(n5287) );
  BUFX2 U798 ( .A(n5661), .Y(n1567) );
  BUFX2 U799 ( .A(n5677), .Y(n1664) );
  BUFX2 U800 ( .A(n5661), .Y(n1568) );
  BUFX2 U801 ( .A(n5671), .Y(n1634) );
  BUFX2 U802 ( .A(n5671), .Y(n1633) );
  BUFX2 U803 ( .A(n5671), .Y(n1632) );
  BUFX2 U804 ( .A(n5671), .Y(n1631) );
  BUFX2 U805 ( .A(n1), .Y(n1563) );
  BUFX2 U806 ( .A(n1), .Y(n1562) );
  BUFX2 U807 ( .A(n1594), .Y(n1581) );
  BUFX2 U808 ( .A(n5663), .Y(n1594) );
  BUFX2 U809 ( .A(n1580), .Y(n1570) );
  BUFX2 U810 ( .A(n1569), .Y(n1580) );
  BUFX2 U811 ( .A(n5661), .Y(n1569) );
  BUFX2 U812 ( .A(n1635), .Y(n1622) );
  BUFX2 U813 ( .A(n5671), .Y(n1635) );
  BUFX2 U814 ( .A(n1677), .Y(n1666) );
  BUFX2 U815 ( .A(n1665), .Y(n1677) );
  BUFX2 U816 ( .A(n5677), .Y(n1665) );
  BUFX2 U817 ( .A(n1), .Y(n1565) );
  BUFX2 U818 ( .A(n1), .Y(n1564) );
  BUFX2 U819 ( .A(n1278), .Y(n1268) );
  BUFX2 U820 ( .A(n1278), .Y(n1266) );
  BUFX2 U821 ( .A(n1278), .Y(n1269) );
  BUFX2 U822 ( .A(n1347), .Y(n1294) );
  BUFX2 U823 ( .A(n1347), .Y(n1293) );
  BUFX2 U824 ( .A(n1348), .Y(n1295) );
  BUFX2 U825 ( .A(n1348), .Y(n1296) );
  BUFX2 U826 ( .A(n1417), .Y(n1351) );
  BUFX2 U827 ( .A(n1418), .Y(n1352) );
  BUFX2 U828 ( .A(n1418), .Y(n1353) );
  BUFX2 U829 ( .A(n1417), .Y(n1350) );
  BUFX2 U830 ( .A(n1418), .Y(n1349) );
  BUFX2 U831 ( .A(n1566), .Y(n1553) );
  BUFX2 U832 ( .A(n1), .Y(n1566) );
  INVX1 U833 ( .A(n1424), .Y(n5760) );
  BUFX2 U834 ( .A(n5757), .Y(n1685) );
  BUFX2 U835 ( .A(n5757), .Y(n1686) );
  BUFX2 U836 ( .A(n5757), .Y(n1689) );
  BUFX2 U837 ( .A(n1292), .Y(n1281) );
  BUFX2 U838 ( .A(n1278), .Y(n1267) );
  BUFX2 U839 ( .A(n1292), .Y(n1280) );
  BUFX2 U840 ( .A(n1292), .Y(n1282) );
  BUFX2 U841 ( .A(n5757), .Y(n1687) );
  BUFX2 U842 ( .A(n5757), .Y(n1688) );
  BUFX2 U843 ( .A(n4005), .Y(n3992) );
  BUFX2 U844 ( .A(n742), .Y(n4005) );
  INVX1 U845 ( .A(n3989), .Y(n3976) );
  NOR2X1 U846 ( .A(n1424), .B(n4597), .Y(n2) );
  INVX1 U847 ( .A(n2), .Y(n5761) );
  BUFX2 U848 ( .A(n1690), .Y(n1678) );
  BUFX2 U849 ( .A(n5757), .Y(n1690) );
  BUFX2 U850 ( .A(n742), .Y(n4004) );
  BUFX2 U851 ( .A(n742), .Y(n4003) );
  BUFX2 U852 ( .A(n742), .Y(n4002) );
  BUFX2 U853 ( .A(n742), .Y(n4001) );
  BUFX2 U854 ( .A(n5759), .Y(n1715) );
  BUFX2 U855 ( .A(n5759), .Y(n1716) );
  BUFX2 U856 ( .A(n5759), .Y(n1713) );
  BUFX2 U857 ( .A(n5759), .Y(n1714) );
  BUFX2 U858 ( .A(n4115), .Y(n4114) );
  BUFX2 U859 ( .A(n736), .Y(n4142) );
  BUFX2 U860 ( .A(n735), .Y(n4170) );
  BUFX2 U861 ( .A(n733), .Y(n4198) );
  BUFX2 U862 ( .A(n729), .Y(n4282) );
  BUFX2 U863 ( .A(n4115), .Y(n4113) );
  BUFX2 U864 ( .A(n736), .Y(n4141) );
  BUFX2 U865 ( .A(n735), .Y(n4169) );
  BUFX2 U866 ( .A(n733), .Y(n4197) );
  BUFX2 U867 ( .A(n4030), .Y(n4028) );
  BUFX2 U868 ( .A(n729), .Y(n4281) );
  BUFX2 U869 ( .A(n727), .Y(n4309) );
  BUFX2 U870 ( .A(n4030), .Y(n4027) );
  BUFX2 U871 ( .A(n739), .Y(n4056) );
  BUFX2 U872 ( .A(n4115), .Y(n4112) );
  BUFX2 U873 ( .A(n736), .Y(n4140) );
  BUFX2 U874 ( .A(n735), .Y(n4168) );
  BUFX2 U875 ( .A(n733), .Y(n4196) );
  BUFX2 U876 ( .A(n729), .Y(n4280) );
  BUFX2 U877 ( .A(n727), .Y(n4308) );
  BUFX2 U878 ( .A(n4059), .Y(n4055) );
  BUFX2 U879 ( .A(n4087), .Y(n4083) );
  BUFX2 U880 ( .A(n4115), .Y(n4111) );
  BUFX2 U881 ( .A(n4143), .Y(n4139) );
  BUFX2 U882 ( .A(n4171), .Y(n4167) );
  BUFX2 U883 ( .A(n4199), .Y(n4195) );
  BUFX2 U884 ( .A(n4283), .Y(n4279) );
  BUFX2 U885 ( .A(n4059), .Y(n4054) );
  BUFX2 U886 ( .A(n4087), .Y(n4082) );
  BUFX2 U887 ( .A(n4115), .Y(n4110) );
  BUFX2 U888 ( .A(n4143), .Y(n4138) );
  BUFX2 U889 ( .A(n4171), .Y(n4166) );
  BUFX2 U890 ( .A(n4199), .Y(n4194) );
  BUFX2 U891 ( .A(n4283), .Y(n4278) );
  BUFX2 U892 ( .A(n4311), .Y(n4306) );
  BUFX2 U893 ( .A(n4059), .Y(n4053) );
  BUFX2 U894 ( .A(n4115), .Y(n4109) );
  BUFX2 U895 ( .A(n4143), .Y(n4137) );
  BUFX2 U896 ( .A(n4171), .Y(n4165) );
  BUFX2 U897 ( .A(n4199), .Y(n4193) );
  BUFX2 U898 ( .A(n4283), .Y(n4277) );
  BUFX2 U899 ( .A(n4311), .Y(n4305) );
  BUFX2 U900 ( .A(n4060), .Y(n4052) );
  BUFX2 U901 ( .A(n4088), .Y(n4080) );
  BUFX2 U902 ( .A(n4116), .Y(n4108) );
  BUFX2 U903 ( .A(n4032), .Y(n4023) );
  BUFX2 U904 ( .A(n4060), .Y(n4051) );
  BUFX2 U905 ( .A(n4088), .Y(n4079) );
  BUFX2 U906 ( .A(n4032), .Y(n4024) );
  BUFX2 U907 ( .A(n4144), .Y(n4136) );
  BUFX2 U908 ( .A(n4172), .Y(n4164) );
  BUFX2 U909 ( .A(n4200), .Y(n4192) );
  BUFX2 U910 ( .A(n4284), .Y(n4276) );
  BUFX2 U911 ( .A(n4312), .Y(n4304) );
  BUFX2 U912 ( .A(n4144), .Y(n4135) );
  BUFX2 U913 ( .A(n4200), .Y(n4191) );
  BUFX2 U914 ( .A(n4284), .Y(n4275) );
  BUFX2 U915 ( .A(n4312), .Y(n4303) );
  BUFX2 U916 ( .A(n4088), .Y(n4078) );
  BUFX2 U917 ( .A(n4116), .Y(n4106) );
  BUFX2 U918 ( .A(n4200), .Y(n4190) );
  BUFX2 U919 ( .A(n4089), .Y(n4077) );
  BUFX2 U920 ( .A(n4145), .Y(n4133) );
  BUFX2 U921 ( .A(n4173), .Y(n4161) );
  BUFX2 U922 ( .A(n4201), .Y(n4189) );
  BUFX2 U923 ( .A(n4285), .Y(n4273) );
  BUFX2 U924 ( .A(n4313), .Y(n4301) );
  BUFX2 U925 ( .A(n4117), .Y(n4104) );
  BUFX2 U926 ( .A(n4285), .Y(n4272) );
  BUFX2 U927 ( .A(n4313), .Y(n4300) );
  BUFX2 U928 ( .A(n4061), .Y(n4047) );
  BUFX2 U929 ( .A(n4117), .Y(n4103) );
  BUFX2 U930 ( .A(n4145), .Y(n4131) );
  BUFX2 U931 ( .A(n4173), .Y(n4159) );
  BUFX2 U932 ( .A(n4201), .Y(n4187) );
  BUFX2 U933 ( .A(n4285), .Y(n4271) );
  BUFX2 U934 ( .A(n3983), .Y(n3988) );
  BUFX2 U935 ( .A(n3984), .Y(n3987) );
  BUFX2 U936 ( .A(n3983), .Y(n3986) );
  BUFX2 U937 ( .A(n3989), .Y(n3985) );
  BUFX2 U938 ( .A(n3989), .Y(n3983) );
  BUFX2 U939 ( .A(n3990), .Y(n3982) );
  BUFX2 U940 ( .A(n3990), .Y(n3981) );
  BUFX2 U941 ( .A(n3990), .Y(n3980) );
  BUFX2 U942 ( .A(n3991), .Y(n3979) );
  BUFX2 U943 ( .A(n3991), .Y(n3978) );
  BUFX2 U944 ( .A(n3991), .Y(n3977) );
  BUFX2 U945 ( .A(n4030), .Y(n4029) );
  BUFX2 U946 ( .A(n4031), .Y(n4026) );
  BUFX2 U947 ( .A(n4311), .Y(n4307) );
  BUFX2 U948 ( .A(n4031), .Y(n4025) );
  BUFX2 U949 ( .A(n4087), .Y(n4081) );
  BUFX2 U950 ( .A(n4116), .Y(n4107) );
  BUFX2 U951 ( .A(n4172), .Y(n4163) );
  BUFX2 U952 ( .A(n4032), .Y(n4022) );
  BUFX2 U953 ( .A(n4060), .Y(n4050) );
  BUFX2 U954 ( .A(n4144), .Y(n4134) );
  BUFX2 U955 ( .A(n4172), .Y(n4162) );
  BUFX2 U956 ( .A(n4284), .Y(n4274) );
  BUFX2 U957 ( .A(n4312), .Y(n4302) );
  BUFX2 U958 ( .A(n4033), .Y(n4021) );
  BUFX2 U959 ( .A(n4061), .Y(n4049) );
  BUFX2 U960 ( .A(n4117), .Y(n4105) );
  BUFX2 U961 ( .A(n4033), .Y(n4020) );
  BUFX2 U962 ( .A(n4061), .Y(n4048) );
  BUFX2 U963 ( .A(n4089), .Y(n4076) );
  BUFX2 U964 ( .A(n4145), .Y(n4132) );
  BUFX2 U965 ( .A(n4173), .Y(n4160) );
  BUFX2 U966 ( .A(n4201), .Y(n4188) );
  BUFX2 U967 ( .A(n4033), .Y(n4019) );
  BUFX2 U968 ( .A(n4089), .Y(n4075) );
  BUFX2 U969 ( .A(n4313), .Y(n4299) );
  BUFX2 U970 ( .A(n3989), .Y(n3984) );
  BUFX2 U971 ( .A(n725), .Y(n4338) );
  BUFX2 U972 ( .A(n4058), .Y(n4057) );
  BUFX2 U973 ( .A(n4087), .Y(n4084) );
  BUFX2 U974 ( .A(n4086), .Y(n4085) );
  BUFX2 U975 ( .A(n725), .Y(n4339) );
  BUFX2 U976 ( .A(n722), .Y(n4367) );
  BUFX2 U977 ( .A(n725), .Y(n4340) );
  BUFX2 U978 ( .A(n722), .Y(n4368) );
  BUFX2 U979 ( .A(n725), .Y(n4341) );
  BUFX2 U980 ( .A(n722), .Y(n4369) );
  INVX1 U981 ( .A(n4031), .Y(n4018) );
  INVX1 U982 ( .A(n4058), .Y(n4046) );
  INVX1 U983 ( .A(n4087), .Y(n4074) );
  INVX1 U984 ( .A(n4108), .Y(n4102) );
  INVX1 U985 ( .A(n4143), .Y(n4130) );
  INVX1 U986 ( .A(n4172), .Y(n4158) );
  INVX1 U987 ( .A(n4199), .Y(n4186) );
  INVX1 U988 ( .A(n4284), .Y(n4270) );
  INVX1 U989 ( .A(n4311), .Y(n4298) );
  BUFX2 U990 ( .A(n730), .Y(n4230) );
  INVX1 U991 ( .A(n4202), .Y(n4229) );
  BUFX2 U992 ( .A(n613), .Y(n1532) );
  BUFX2 U993 ( .A(n701), .Y(n1444) );
  BUFX2 U994 ( .A(n669), .Y(n1476) );
  BUFX2 U995 ( .A(n637), .Y(n1508) );
  BUFX2 U996 ( .A(n709), .Y(n1436) );
  BUFX2 U997 ( .A(n677), .Y(n1468) );
  BUFX2 U998 ( .A(n645), .Y(n1500) );
  XOR2XL U999 ( .A(n4819), .B(new_sboxw[6]), .Y(n4820) );
  XOR2XL U1000 ( .A(n4807), .B(new_sboxw[6]), .Y(n4808) );
  XOR2XL U1001 ( .A(n4818), .B(new_sboxw[6]), .Y(n4800) );
  XOR2XL U1002 ( .A(n5081), .B(new_sboxw[6]), .Y(n5713) );
  XOR2XL U1003 ( .A(n5069), .B(new_sboxw[6]), .Y(n5714) );
  XOR2XL U1004 ( .A(n4884), .B(new_sboxw[0]), .Y(n5730) );
  XOR2XL U1005 ( .A(n4872), .B(new_sboxw[0]), .Y(n5731) );
  OAI221XL U1006 ( .A0(n941), .A1(n3995), .B0(n3942), .B1(n5865), .C0(n942), 
        .Y(n642) );
  INVX1 U1007 ( .A(n1420), .Y(n942) );
  OAI222XL U1008 ( .A0(n4598), .A1(n1421), .B0(n5066), .B1(n5678), .C0(n4593), 
        .C1(n4), .Y(n1420) );
  BUFX2 U1009 ( .A(n648), .Y(n1497) );
  BUFX2 U1010 ( .A(n680), .Y(n1465) );
  BUFX2 U1011 ( .A(n674), .Y(n1471) );
  INVX1 U1012 ( .A(n5079), .Y(n1071) );
  BUFX2 U1013 ( .A(n714), .Y(n1431) );
  BUFX2 U1014 ( .A(n712), .Y(n1433) );
  BUFX2 U1015 ( .A(n706), .Y(n1439) );
  BUFX2 U1016 ( .A(n688), .Y(n1457) );
  BUFX2 U1017 ( .A(n682), .Y(n1463) );
  BUFX2 U1018 ( .A(n656), .Y(n1489) );
  BUFX2 U1019 ( .A(n650), .Y(n1495) );
  BUFX2 U1020 ( .A(n624), .Y(n1521) );
  BUFX2 U1021 ( .A(n610), .Y(n1535) );
  BUFX2 U1022 ( .A(n605), .Y(n1540) );
  INVX1 U1023 ( .A(n8), .Y(n1421) );
  INVX1 U1024 ( .A(n5068), .Y(n815) );
  INVX1 U1025 ( .A(n4871), .Y(n839) );
  INVX1 U1026 ( .A(n4882), .Y(n1095) );
  INVX1 U1027 ( .A(n5112), .Y(n1067) );
  BUFX2 U1028 ( .A(n720), .Y(n1425) );
  BUFX2 U1029 ( .A(n705), .Y(n1440) );
  BUFX2 U1030 ( .A(n699), .Y(n1446) );
  BUFX2 U1031 ( .A(n697), .Y(n1448) );
  BUFX2 U1032 ( .A(n673), .Y(n1472) );
  BUFX2 U1033 ( .A(n618), .Y(n1527) );
  BUFX2 U1034 ( .A(n616), .Y(n1529) );
  XOR2XL U1035 ( .A(n4692), .B(new_sboxw[2]), .Y(n4693) );
  XOR2XL U1036 ( .A(n4724), .B(new_sboxw[3]), .Y(n4725) );
  XOR2XL U1037 ( .A(n4788), .B(new_sboxw[5]), .Y(n4789) );
  XOR2XL U1038 ( .A(n4851), .B(new_sboxw[7]), .Y(n4852) );
  XOR2XL U1039 ( .A(n4950), .B(new_sboxw[10]), .Y(n4951) );
  XOR2XL U1040 ( .A(n5049), .B(new_sboxw[13]), .Y(n5050) );
  XOR2XL U1041 ( .A(n5114), .B(new_sboxw[15]), .Y(n5115) );
  XOR2XL U1042 ( .A(n4680), .B(new_sboxw[2]), .Y(n4681) );
  XOR2XL U1043 ( .A(n4712), .B(new_sboxw[3]), .Y(n4713) );
  XOR2XL U1044 ( .A(n4776), .B(new_sboxw[5]), .Y(n4777) );
  XOR2XL U1045 ( .A(n4839), .B(new_sboxw[7]), .Y(n4840) );
  XOR2XL U1046 ( .A(n4938), .B(new_sboxw[10]), .Y(n4939) );
  XOR2XL U1047 ( .A(n5037), .B(new_sboxw[13]), .Y(n5038) );
  XOR2XL U1048 ( .A(n5102), .B(new_sboxw[15]), .Y(n5103) );
  XOR2XL U1049 ( .A(n4691), .B(new_sboxw[2]), .Y(n4673) );
  XOR2XL U1050 ( .A(n4723), .B(new_sboxw[3]), .Y(n4705) );
  XOR2XL U1051 ( .A(n4787), .B(new_sboxw[5]), .Y(n4769) );
  XOR2XL U1052 ( .A(n4850), .B(new_sboxw[7]), .Y(n4832) );
  XOR2XL U1053 ( .A(n4949), .B(new_sboxw[10]), .Y(n4931) );
  XOR2XL U1054 ( .A(n5048), .B(new_sboxw[13]), .Y(n5030) );
  XOR2XL U1055 ( .A(n5113), .B(new_sboxw[15]), .Y(n5095) );
  XOR2XL U1056 ( .A(n4917), .B(new_sboxw[9]), .Y(n4918) );
  XOR2XL U1057 ( .A(n4905), .B(new_sboxw[9]), .Y(n4906) );
  XOR2XL U1058 ( .A(n4916), .B(new_sboxw[9]), .Y(n4898) );
  XOR2XL U1059 ( .A(n4950), .B(new_sboxw[2]), .Y(n5724) );
  XOR2XL U1060 ( .A(n4983), .B(new_sboxw[3]), .Y(n5721) );
  XOR2XL U1061 ( .A(n5049), .B(new_sboxw[5]), .Y(n5715) );
  XOR2XL U1062 ( .A(n5114), .B(new_sboxw[7]), .Y(n5710) );
  XOR2XL U1063 ( .A(n5213), .B(new_sboxw[10]), .Y(n5701) );
  XOR2XL U1064 ( .A(n5312), .B(new_sboxw[13]), .Y(n5692) );
  XOR2XL U1065 ( .A(n5377), .B(new_sboxw[15]), .Y(n5687) );
  XOR2XL U1066 ( .A(n4938), .B(new_sboxw[2]), .Y(n5725) );
  XOR2XL U1067 ( .A(n4971), .B(new_sboxw[3]), .Y(n5722) );
  XOR2XL U1068 ( .A(n5037), .B(new_sboxw[5]), .Y(n5716) );
  XOR2XL U1069 ( .A(n5102), .B(new_sboxw[7]), .Y(n5711) );
  XOR2XL U1070 ( .A(n5201), .B(new_sboxw[10]), .Y(n5702) );
  XOR2XL U1071 ( .A(n5300), .B(new_sboxw[13]), .Y(n5693) );
  XOR2XL U1072 ( .A(n5365), .B(new_sboxw[15]), .Y(n5688) );
  XOR2XL U1073 ( .A(n4949), .B(new_sboxw[2]), .Y(n5726) );
  XOR2XL U1074 ( .A(n4982), .B(new_sboxw[3]), .Y(n5723) );
  XOR2XL U1075 ( .A(n5048), .B(new_sboxw[5]), .Y(n5717) );
  XOR2XL U1076 ( .A(n5113), .B(new_sboxw[7]), .Y(n5712) );
  XOR2XL U1077 ( .A(n5212), .B(new_sboxw[10]), .Y(n5703) );
  XOR2XL U1078 ( .A(n5311), .B(new_sboxw[13]), .Y(n5694) );
  XOR2XL U1079 ( .A(n5376), .B(new_sboxw[15]), .Y(n5689) );
  XOR2XL U1080 ( .A(n5180), .B(new_sboxw[9]), .Y(n5704) );
  XOR2XL U1081 ( .A(n5081), .B(new_sboxw[14]), .Y(n5082) );
  XOR2XL U1082 ( .A(n5069), .B(new_sboxw[14]), .Y(n5070) );
  XOR2XL U1083 ( .A(n5343), .B(new_sboxw[14]), .Y(n5691) );
  XOR2XL U1084 ( .A(n5179), .B(new_sboxw[9]), .Y(n5706) );
  XOR2X1 U1085 ( .A(n4756), .B(new_sboxw[28]), .Y(n5742) );
  XOR2X1 U1086 ( .A(n4744), .B(new_sboxw[28]), .Y(n5743) );
  XOR2X1 U1087 ( .A(n4755), .B(new_sboxw[28]), .Y(n5744) );
  XOR2X1 U1088 ( .A(n4819), .B(new_sboxw[30]), .Y(n5736) );
  XOR2X1 U1089 ( .A(n4807), .B(new_sboxw[30]), .Y(n5737) );
  XOR2X1 U1090 ( .A(n4818), .B(new_sboxw[30]), .Y(n5738) );
  XOR2X1 U1091 ( .A(n4628), .B(new_sboxw[24]), .Y(n5754) );
  XOR2X1 U1092 ( .A(n4660), .B(new_sboxw[25]), .Y(n5751) );
  XOR2X1 U1093 ( .A(n4617), .B(new_sboxw[24]), .Y(n5755) );
  XOR2X1 U1094 ( .A(n4648), .B(new_sboxw[25]), .Y(n5752) );
  XOR2X1 U1095 ( .A(n4627), .B(new_sboxw[24]), .Y(n5756) );
  XOR2X1 U1096 ( .A(n4659), .B(new_sboxw[25]), .Y(n5753) );
  XOR2XL U1097 ( .A(n5267), .B(new_sboxw[12]), .Y(n5696) );
  XOR2XL U1098 ( .A(n5147), .B(new_sboxw[8]), .Y(n5707) );
  XOR2XL U1099 ( .A(n5135), .B(new_sboxw[8]), .Y(n5708) );
  XOR2XL U1100 ( .A(n4905), .B(new_sboxw[1]), .Y(n5728) );
  XOR2XL U1101 ( .A(n4916), .B(new_sboxw[1]), .Y(n5729) );
  XOR2XL U1102 ( .A(n4660), .B(new_sboxw[1]), .Y(n4661) );
  XOR2XL U1103 ( .A(n4648), .B(new_sboxw[1]), .Y(n4649) );
  XOR2XL U1104 ( .A(n4659), .B(new_sboxw[1]), .Y(n4641) );
  XOR2XL U1105 ( .A(n5146), .B(new_sboxw[8]), .Y(n5709) );
  XOR2XL U1106 ( .A(n4864), .B(new_sboxw[8]), .Y(n837) );
  XOR2XL U1107 ( .A(n4883), .B(new_sboxw[8]), .Y(n4865) );
  XOR2X1 U1108 ( .A(n4724), .B(new_sboxw[27]), .Y(n5745) );
  XOR2X1 U1109 ( .A(n4788), .B(new_sboxw[29]), .Y(n5739) );
  XOR2X1 U1110 ( .A(n4851), .B(new_sboxw[31]), .Y(n5733) );
  XOR2X1 U1111 ( .A(n4712), .B(new_sboxw[27]), .Y(n5746) );
  XOR2X1 U1112 ( .A(n4776), .B(new_sboxw[29]), .Y(n5740) );
  XOR2X1 U1113 ( .A(n4839), .B(new_sboxw[31]), .Y(n5734) );
  XOR2X1 U1114 ( .A(n4723), .B(new_sboxw[27]), .Y(n5747) );
  XOR2X1 U1115 ( .A(n4787), .B(new_sboxw[29]), .Y(n5741) );
  XOR2X1 U1116 ( .A(n4850), .B(new_sboxw[31]), .Y(n5735) );
  XOR2X1 U1117 ( .A(n5666), .B(new_sboxw[31]), .Y(n1129) );
  XOR2X1 U1118 ( .A(n5652), .B(new_sboxw[31]), .Y(n1001) );
  XOR2X1 U1119 ( .A(n5664), .B(new_sboxw[31]), .Y(n873) );
  XOR2X1 U1120 ( .A(n5434), .B(n5435), .Y(n5448) );
  XOR2X1 U1121 ( .A(n5542), .B(n5543), .Y(n5556) );
  XOR2X1 U1122 ( .A(n5578), .B(n5579), .Y(n5592) );
  XOR2X1 U1123 ( .A(n5614), .B(n5615), .Y(n5628) );
  XOR2X1 U1124 ( .A(n5506), .B(n5507), .Y(n5520) );
  XOR2X1 U1125 ( .A(n5470), .B(n5471), .Y(n5484) );
  XOR2X1 U1126 ( .A(n5398), .B(n5399), .Y(n5412) );
  XOR2X1 U1127 ( .A(n5377), .B(new_sboxw[23]), .Y(n5378) );
  XOR2X1 U1128 ( .A(n5365), .B(new_sboxw[23]), .Y(n5366) );
  XOR2X1 U1129 ( .A(n5376), .B(new_sboxw[23]), .Y(n5358) );
  XOR2X1 U1130 ( .A(n5357), .B(new_sboxw[23]), .Y(n777) );
  XOR2X1 U1131 ( .A(n5666), .B(n5665), .Y(n5679) );
  XOR2X1 U1132 ( .A(n5652), .B(n5665), .Y(n5681) );
  XOR2X1 U1133 ( .A(n5664), .B(n5665), .Y(n5683) );
  XNOR2X1 U1134 ( .A(n5447), .B(n5446), .Y(n5430) );
  XNOR2X1 U1135 ( .A(n5555), .B(n5554), .Y(n5538) );
  XNOR2X1 U1136 ( .A(n5591), .B(n5590), .Y(n5574) );
  XNOR2X1 U1137 ( .A(n5627), .B(n5626), .Y(n5610) );
  XNOR2X1 U1138 ( .A(n5519), .B(n5518), .Y(n5502) );
  XNOR2X1 U1139 ( .A(n5483), .B(n5482), .Y(n5466) );
  XNOR2X1 U1140 ( .A(n5411), .B(n5410), .Y(n5394) );
  XNOR2X1 U1141 ( .A(n5447), .B(n5436), .Y(n5440) );
  XNOR2X1 U1142 ( .A(n5555), .B(n5544), .Y(n5548) );
  XNOR2X1 U1143 ( .A(n5591), .B(n5580), .Y(n5584) );
  XNOR2X1 U1144 ( .A(n5627), .B(n5616), .Y(n5620) );
  XNOR2X1 U1145 ( .A(n5519), .B(n5508), .Y(n5512) );
  XNOR2X1 U1146 ( .A(n5483), .B(n5472), .Y(n5476) );
  XNOR2X1 U1147 ( .A(n5411), .B(n5400), .Y(n5404) );
  XNOR2X1 U1148 ( .A(n5447), .B(n5449), .Y(n5453) );
  XNOR2X1 U1149 ( .A(n5555), .B(n5557), .Y(n5561) );
  XNOR2X1 U1150 ( .A(n5591), .B(n5593), .Y(n5597) );
  XNOR2X1 U1151 ( .A(n5627), .B(n5629), .Y(n5633) );
  XNOR2X1 U1152 ( .A(n5519), .B(n5521), .Y(n5525) );
  XNOR2X1 U1153 ( .A(n5483), .B(n5485), .Y(n5489) );
  XNOR2X1 U1154 ( .A(n5411), .B(n5413), .Y(n5417) );
  XOR2X1 U1155 ( .A(n5651), .B(n5665), .Y(n5684) );
  BUFX2 U1156 ( .A(n672), .Y(n1473) );
  BUFX2 U1157 ( .A(n711), .Y(n1434) );
  BUFX2 U1158 ( .A(n679), .Y(n1466) );
  BUFX2 U1159 ( .A(n676), .Y(n1469) );
  BUFX2 U1160 ( .A(n668), .Y(n1477) );
  BUFX2 U1161 ( .A(n647), .Y(n1498) );
  BUFX2 U1162 ( .A(n644), .Y(n1501) );
  INVX1 U1163 ( .A(n5642), .Y(n5665) );
  BUFX2 U1164 ( .A(n703), .Y(n1442) );
  BUFX2 U1165 ( .A(n704), .Y(n1441) );
  INVX1 U1166 ( .A(n5411), .Y(n5399) );
  INVX1 U1167 ( .A(n5519), .Y(n5507) );
  INVX1 U1168 ( .A(n5483), .Y(n5471) );
  INVX1 U1169 ( .A(n5447), .Y(n5435) );
  INVX1 U1170 ( .A(n5555), .Y(n5543) );
  INVX1 U1171 ( .A(n5591), .Y(n5579) );
  INVX1 U1172 ( .A(n5627), .Y(n5615) );
  INVX1 U1173 ( .A(n4904), .Y(n835) );
  BUFX2 U1174 ( .A(n708), .Y(n1437) );
  BUFX2 U1175 ( .A(n640), .Y(n1505) );
  BUFX2 U1176 ( .A(n700), .Y(n1445) );
  BUFX2 U1177 ( .A(n634), .Y(n1511) );
  OAI221XL U1178 ( .A0(n1037), .A1(n3993), .B0(n3940), .B1(n5873), .C0(n1038), 
        .Y(n666) );
  INVX1 U1179 ( .A(n5334), .Y(n1037) );
  INVX1 U1180 ( .A(n1423), .Y(n1038) );
  OAI222XL U1181 ( .A0(n4598), .A1(n5342), .B0(n5337), .B1(n5678), .C0(n4593), 
        .C1(n5), .Y(n1423) );
  INVX1 U1182 ( .A(n5003), .Y(n823) );
  INVX1 U1183 ( .A(n4775), .Y(n851) );
  INVX1 U1184 ( .A(n4806), .Y(n847) );
  INVX1 U1185 ( .A(n4838), .Y(n843) );
  INVX1 U1186 ( .A(n4937), .Y(n831) );
  INVX1 U1187 ( .A(n4970), .Y(n827) );
  INVX1 U1188 ( .A(n5036), .Y(n819) );
  INVX1 U1189 ( .A(n4743), .Y(n855) );
  INVX1 U1190 ( .A(n5101), .Y(n811) );
  INVX1 U1191 ( .A(n5134), .Y(n807) );
  INVX1 U1192 ( .A(n5167), .Y(n803) );
  INVX1 U1193 ( .A(n5200), .Y(n799) );
  INVX1 U1194 ( .A(n5266), .Y(n791) );
  INVX1 U1195 ( .A(n5299), .Y(n787) );
  INVX1 U1196 ( .A(n5332), .Y(n783) );
  INVX1 U1197 ( .A(n5364), .Y(n779) );
  BUFX2 U1198 ( .A(n671), .Y(n1474) );
  INVX1 U1199 ( .A(n4690), .Y(n1119) );
  INVX1 U1200 ( .A(n4722), .Y(n1115) );
  INVX1 U1201 ( .A(n4754), .Y(n1111) );
  INVX1 U1202 ( .A(n4786), .Y(n1107) );
  INVX1 U1203 ( .A(n4817), .Y(n1103) );
  INVX1 U1204 ( .A(n4849), .Y(n1099) );
  INVX1 U1205 ( .A(n4948), .Y(n1087) );
  INVX1 U1206 ( .A(n4981), .Y(n1083) );
  INVX1 U1207 ( .A(n5047), .Y(n1075) );
  INVX1 U1208 ( .A(n5211), .Y(n1055) );
  INVX1 U1209 ( .A(n5310), .Y(n1043) );
  INVX1 U1210 ( .A(n5375), .Y(n1035) );
  INVX1 U1211 ( .A(n4626), .Y(n1127) );
  INVX1 U1212 ( .A(n4658), .Y(n1123) );
  INVX1 U1213 ( .A(n4915), .Y(n1091) );
  INVX1 U1214 ( .A(n5145), .Y(n1063) );
  INVX1 U1215 ( .A(n5178), .Y(n1059) );
  INVX1 U1216 ( .A(n5277), .Y(n1047) );
  INVX1 U1217 ( .A(n5014), .Y(n1079) );
  BUFX2 U1218 ( .A(n695), .Y(n1450) );
  BUFX2 U1219 ( .A(n663), .Y(n1482) );
  BUFX2 U1220 ( .A(n631), .Y(n1514) );
  BUFX2 U1221 ( .A(n599), .Y(n1546) );
  BUFX2 U1222 ( .A(n692), .Y(n1453) );
  BUFX2 U1223 ( .A(n660), .Y(n1485) );
  BUFX2 U1224 ( .A(n628), .Y(n1517) );
  BUFX2 U1225 ( .A(n596), .Y(n1549) );
  BUFX2 U1226 ( .A(n691), .Y(n1454) );
  BUFX2 U1227 ( .A(n659), .Y(n1486) );
  BUFX2 U1228 ( .A(n627), .Y(n1518) );
  BUFX2 U1229 ( .A(n595), .Y(n1550) );
  BUFX2 U1230 ( .A(n690), .Y(n1455) );
  BUFX2 U1231 ( .A(n658), .Y(n1487) );
  BUFX2 U1232 ( .A(n626), .Y(n1519) );
  BUFX2 U1233 ( .A(n594), .Y(n1551) );
  BUFX2 U1234 ( .A(n693), .Y(n1452) );
  BUFX2 U1235 ( .A(n661), .Y(n1484) );
  BUFX2 U1236 ( .A(n629), .Y(n1516) );
  BUFX2 U1237 ( .A(n597), .Y(n1548) );
  BUFX2 U1238 ( .A(n694), .Y(n1451) );
  BUFX2 U1239 ( .A(n662), .Y(n1483) );
  BUFX2 U1240 ( .A(n630), .Y(n1515) );
  BUFX2 U1241 ( .A(n598), .Y(n1547) );
  BUFX2 U1242 ( .A(n696), .Y(n1449) );
  BUFX2 U1243 ( .A(n664), .Y(n1481) );
  BUFX2 U1244 ( .A(n632), .Y(n1513) );
  BUFX2 U1245 ( .A(n600), .Y(n1545) );
  BUFX2 U1246 ( .A(n689), .Y(n1456) );
  BUFX2 U1247 ( .A(n657), .Y(n1488) );
  BUFX2 U1248 ( .A(n625), .Y(n1520) );
  BUFX2 U1249 ( .A(n593), .Y(n1552) );
  BUFX2 U1250 ( .A(n719), .Y(n1426) );
  BUFX2 U1251 ( .A(n718), .Y(n1427) );
  BUFX2 U1252 ( .A(n717), .Y(n1428) );
  BUFX2 U1253 ( .A(n715), .Y(n1430) );
  BUFX2 U1254 ( .A(n713), .Y(n1432) );
  BUFX2 U1255 ( .A(n710), .Y(n1435) );
  BUFX2 U1256 ( .A(n707), .Y(n1438) );
  BUFX2 U1257 ( .A(n702), .Y(n1443) );
  BUFX2 U1258 ( .A(n698), .Y(n1447) );
  BUFX2 U1259 ( .A(n687), .Y(n1458) );
  BUFX2 U1260 ( .A(n686), .Y(n1459) );
  BUFX2 U1261 ( .A(n685), .Y(n1460) );
  BUFX2 U1262 ( .A(n684), .Y(n1461) );
  BUFX2 U1263 ( .A(n683), .Y(n1462) );
  BUFX2 U1264 ( .A(n681), .Y(n1464) );
  BUFX2 U1265 ( .A(n678), .Y(n1467) );
  BUFX2 U1266 ( .A(n675), .Y(n1470) );
  BUFX2 U1267 ( .A(n670), .Y(n1475) );
  BUFX2 U1268 ( .A(n667), .Y(n1478) );
  BUFX2 U1269 ( .A(n665), .Y(n1480) );
  BUFX2 U1270 ( .A(n655), .Y(n1490) );
  BUFX2 U1271 ( .A(n654), .Y(n1491) );
  BUFX2 U1272 ( .A(n653), .Y(n1492) );
  BUFX2 U1273 ( .A(n652), .Y(n1493) );
  BUFX2 U1274 ( .A(n651), .Y(n1494) );
  BUFX2 U1275 ( .A(n649), .Y(n1496) );
  BUFX2 U1276 ( .A(n646), .Y(n1499) );
  BUFX2 U1277 ( .A(n643), .Y(n1502) );
  BUFX2 U1278 ( .A(n641), .Y(n1504) );
  BUFX2 U1279 ( .A(n639), .Y(n1506) );
  BUFX2 U1280 ( .A(n638), .Y(n1507) );
  BUFX2 U1281 ( .A(n636), .Y(n1509) );
  BUFX2 U1282 ( .A(n635), .Y(n1510) );
  BUFX2 U1283 ( .A(n633), .Y(n1512) );
  BUFX2 U1284 ( .A(n623), .Y(n1522) );
  BUFX2 U1285 ( .A(n622), .Y(n1523) );
  BUFX2 U1286 ( .A(n621), .Y(n1524) );
  BUFX2 U1287 ( .A(n620), .Y(n1525) );
  BUFX2 U1288 ( .A(n619), .Y(n1526) );
  BUFX2 U1289 ( .A(n617), .Y(n1528) );
  BUFX2 U1290 ( .A(n615), .Y(n1530) );
  BUFX2 U1291 ( .A(n614), .Y(n1531) );
  BUFX2 U1292 ( .A(n612), .Y(n1533) );
  BUFX2 U1293 ( .A(n611), .Y(n1534) );
  BUFX2 U1294 ( .A(n609), .Y(n1536) );
  BUFX2 U1295 ( .A(n608), .Y(n1537) );
  BUFX2 U1296 ( .A(n607), .Y(n1538) );
  BUFX2 U1297 ( .A(n606), .Y(n1539) );
  BUFX2 U1298 ( .A(n604), .Y(n1541) );
  BUFX2 U1299 ( .A(n603), .Y(n1542) );
  BUFX2 U1300 ( .A(n602), .Y(n1543) );
  BUFX2 U1301 ( .A(n601), .Y(n1544) );
  BUFX2 U1302 ( .A(n716), .Y(n1429) );
  XOR2X1 U1303 ( .A(n5557), .B(new_sboxw[28]), .Y(n1141) );
  XOR2X1 U1304 ( .A(n5544), .B(new_sboxw[28]), .Y(n1013) );
  XOR2X1 U1305 ( .A(n5554), .B(new_sboxw[28]), .Y(n885) );
  XOR2XL U1306 ( .A(n4744), .B(new_sboxw[4]), .Y(n4745) );
  XOR2X1 U1307 ( .A(n5629), .B(new_sboxw[30]), .Y(n1133) );
  XOR2X1 U1308 ( .A(n5616), .B(new_sboxw[30]), .Y(n1005) );
  XOR2X1 U1309 ( .A(n5626), .B(new_sboxw[30]), .Y(n877) );
  XOR2X1 U1310 ( .A(n5449), .B(new_sboxw[25]), .Y(n1153) );
  XOR2X1 U1311 ( .A(n5436), .B(new_sboxw[25]), .Y(n1025) );
  XOR2X1 U1312 ( .A(n5446), .B(new_sboxw[25]), .Y(n897) );
  XOR2X1 U1313 ( .A(n5413), .B(new_sboxw[24]), .Y(n1157) );
  XOR2X1 U1314 ( .A(n5400), .B(new_sboxw[24]), .Y(n1029) );
  XOR2X1 U1315 ( .A(n5410), .B(new_sboxw[24]), .Y(n901) );
  XOR2XL U1316 ( .A(n5278), .B(new_sboxw[12]), .Y(n5697) );
  XOR2X1 U1317 ( .A(n5279), .B(new_sboxw[20]), .Y(n5280) );
  XOR2X1 U1318 ( .A(n5267), .B(new_sboxw[20]), .Y(n5268) );
  XOR2X1 U1319 ( .A(n5278), .B(new_sboxw[20]), .Y(n5260) );
  XOR2XL U1320 ( .A(n5016), .B(new_sboxw[4]), .Y(n5718) );
  XOR2X1 U1321 ( .A(n5259), .B(new_sboxw[20]), .Y(n789) );
  XOR2XL U1322 ( .A(n5004), .B(new_sboxw[4]), .Y(n5719) );
  XOR2XL U1323 ( .A(n5015), .B(new_sboxw[4]), .Y(n5720) );
  XOR2XL U1324 ( .A(n4736), .B(new_sboxw[4]), .Y(n853) );
  XOR2X1 U1325 ( .A(n5344), .B(new_sboxw[22]), .Y(n5345) );
  XOR2X1 U1326 ( .A(n5333), .B(new_sboxw[22]), .Y(n5334) );
  XOR2X1 U1327 ( .A(n5343), .B(new_sboxw[22]), .Y(n5326) );
  XOR2X1 U1328 ( .A(n5135), .B(new_sboxw[16]), .Y(n5136) );
  XOR2X1 U1329 ( .A(n5147), .B(new_sboxw[16]), .Y(n5148) );
  XOR2X1 U1330 ( .A(n5180), .B(new_sboxw[17]), .Y(n5181) );
  XOR2X1 U1331 ( .A(n5168), .B(new_sboxw[17]), .Y(n5169) );
  XOR2X1 U1332 ( .A(n5146), .B(new_sboxw[16]), .Y(n5128) );
  XOR2X1 U1333 ( .A(n5179), .B(new_sboxw[17]), .Y(n5161) );
  XOR2X1 U1334 ( .A(n5325), .B(new_sboxw[22]), .Y(n781) );
  XOR2X1 U1335 ( .A(n5127), .B(new_sboxw[16]), .Y(n805) );
  XOR2X1 U1336 ( .A(n5160), .B(new_sboxw[17]), .Y(n801) );
  XOR2X1 U1337 ( .A(n4692), .B(new_sboxw[26]), .Y(n5748) );
  XOR2X1 U1338 ( .A(n4680), .B(new_sboxw[26]), .Y(n5749) );
  XOR2X1 U1339 ( .A(n4691), .B(new_sboxw[26]), .Y(n5750) );
  XOR2X1 U1340 ( .A(n5593), .B(new_sboxw[29]), .Y(n1137) );
  XOR2X1 U1341 ( .A(n5580), .B(new_sboxw[29]), .Y(n1009) );
  XOR2X1 U1342 ( .A(n5590), .B(new_sboxw[29]), .Y(n881) );
  XOR2X1 U1343 ( .A(n5521), .B(new_sboxw[27]), .Y(n1145) );
  XOR2X1 U1344 ( .A(n5508), .B(new_sboxw[27]), .Y(n1017) );
  XOR2X1 U1345 ( .A(n5518), .B(new_sboxw[27]), .Y(n889) );
  XOR2X1 U1346 ( .A(n5485), .B(new_sboxw[26]), .Y(n1149) );
  XOR2X1 U1347 ( .A(n5472), .B(new_sboxw[26]), .Y(n1021) );
  XOR2X1 U1348 ( .A(n5482), .B(new_sboxw[26]), .Y(n893) );
  XOR2X1 U1349 ( .A(n5213), .B(new_sboxw[18]), .Y(n5214) );
  XOR2X1 U1350 ( .A(n5246), .B(new_sboxw[19]), .Y(n5247) );
  XOR2X1 U1351 ( .A(n5312), .B(new_sboxw[21]), .Y(n5313) );
  XOR2X1 U1352 ( .A(n5201), .B(new_sboxw[18]), .Y(n5202) );
  XOR2X1 U1353 ( .A(n5234), .B(new_sboxw[19]), .Y(n5235) );
  XOR2X1 U1354 ( .A(n5300), .B(new_sboxw[21]), .Y(n5301) );
  XOR2X1 U1355 ( .A(n5212), .B(new_sboxw[18]), .Y(n5194) );
  XOR2X1 U1356 ( .A(n5245), .B(new_sboxw[19]), .Y(n5227) );
  XOR2X1 U1357 ( .A(n5311), .B(new_sboxw[21]), .Y(n5293) );
  XOR2X1 U1358 ( .A(n5193), .B(new_sboxw[18]), .Y(n797) );
  XOR2X1 U1359 ( .A(n5226), .B(new_sboxw[19]), .Y(n793) );
  XOR2X1 U1360 ( .A(n5292), .B(new_sboxw[21]), .Y(n785) );
  NAND2BX1 U1361 ( .AN(n5678), .B(n4425), .Y(n5677) );
  NAND2BX1 U1362 ( .AN(n4591), .B(n4435), .Y(n5661) );
  NAND3BX1 U1363 ( .AN(n3934), .B(n4600), .C(n4436), .Y(n4601) );
  INVX1 U1364 ( .A(n4616), .Y(n871) );
  INVX1 U1365 ( .A(n4679), .Y(n863) );
  INVX1 U1366 ( .A(n4711), .Y(n859) );
  INVX1 U1367 ( .A(n4647), .Y(n867) );
  INVX1 U1368 ( .A(n769), .Y(n5420) );
  INVX1 U1369 ( .A(n757), .Y(n5528) );
  INVX1 U1370 ( .A(n753), .Y(n5564) );
  INVX1 U1371 ( .A(n749), .Y(n5600) );
  INVX1 U1372 ( .A(n761), .Y(n5492) );
  INVX1 U1373 ( .A(n765), .Y(n5456) );
  INVX1 U1374 ( .A(n773), .Y(n5384) );
  OAI222XL U1375 ( .A0(n5768), .A1(n1587), .B0(n1575), .B1(n5426), .C0(n1555), 
        .C1(n5425), .Y(n3664) );
  OAI222XL U1376 ( .A0(n5830), .A1(n1588), .B0(n1574), .B1(n5534), .C0(n1554), 
        .C1(n5533), .Y(n3661) );
  OAI222XL U1377 ( .A0(n5846), .A1(n1588), .B0(n1573), .B1(n5570), .C0(n1554), 
        .C1(n5569), .Y(n3660) );
  OAI222XL U1378 ( .A0(n5862), .A1(n1589), .B0(n1573), .B1(n5606), .C0(n1553), 
        .C1(n5605), .Y(n3659) );
  OAI222XL U1379 ( .A0(n5814), .A1(n1587), .B0(n1574), .B1(n5498), .C0(n1554), 
        .C1(n5497), .Y(n3662) );
  OAI222XL U1380 ( .A0(n5798), .A1(n1587), .B0(n1574), .B1(n5462), .C0(n1555), 
        .C1(n5461), .Y(n3663) );
  OAI222XL U1381 ( .A0(n5782), .A1(n1586), .B0(n1575), .B1(n5390), .C0(n1564), 
        .C1(n5389), .Y(n3665) );
  OAI222XL U1382 ( .A0(n5878), .A1(n1589), .B0(n1573), .B1(n5643), .C0(n1553), 
        .C1(n5641), .Y(n3658) );
  BUFX2 U1383 ( .A(N32), .Y(n1347) );
  BUFX2 U1384 ( .A(N32), .Y(n1348) );
  BUFX2 U1385 ( .A(N34), .Y(n1278) );
  BUFX2 U1386 ( .A(N31), .Y(n1417) );
  BUFX2 U1387 ( .A(N31), .Y(n1418) );
  BUFX2 U1388 ( .A(n1265), .Y(n1276) );
  BUFX2 U1389 ( .A(n1277), .Y(n1265) );
  BUFX2 U1390 ( .A(N34), .Y(n1277) );
  AO21X1 U1391 ( .A0(n279), .A1(round_ctr_reg[0]), .B0(n4588), .Y(n4594) );
  NAND2BX1 U1392 ( .AN(round_ctr_reg[0]), .B(n1721), .Y(n4597) );
  INVX1 U1393 ( .A(n4591), .Y(n4592) );
  BUFX2 U1394 ( .A(n5763), .Y(n1424) );
  BUFX2 U1395 ( .A(N33), .Y(n1291) );
  BUFX2 U1396 ( .A(N33), .Y(n1292) );
  INVX1 U1397 ( .A(n1721), .Y(n4588) );
  BUFX2 U1398 ( .A(n1279), .Y(n1289) );
  BUFX2 U1399 ( .A(n1290), .Y(n1279) );
  BUFX2 U1400 ( .A(N33), .Y(n1290) );
  INVX1 U1401 ( .A(n4600), .Y(n4602) );
  NAND2X1 U1402 ( .A(n5760), .B(n1723), .Y(n1722) );
  NAND2X1 U1403 ( .A(n1722), .B(n1723), .Y(n1726) );
  NAND2X1 U1404 ( .A(n723), .B(n724), .Y(n722) );
  NAND2BX1 U1405 ( .AN(n731), .B(n723), .Y(n730) );
  NAND2X1 U1406 ( .A(n726), .B(n724), .Y(n725) );
  NAND2X1 U1407 ( .A(n5763), .B(n1733), .Y(n1732) );
  BUFX2 U1408 ( .A(n727), .Y(n4310) );
  INVX1 U1409 ( .A(n5764), .Y(n734) );
  BUFX2 U1410 ( .A(n739), .Y(n4058) );
  BUFX2 U1411 ( .A(n732), .Y(n4202) );
  NOR2BX1 U1412 ( .AN(n726), .B(n731), .Y(n732) );
  BUFX2 U1413 ( .A(n5762), .Y(n3989) );
  BUFX2 U1414 ( .A(n5762), .Y(n3990) );
  BUFX2 U1415 ( .A(n5762), .Y(n3991) );
  AO22X1 U1416 ( .A0(n5760), .A1(n279), .B0(n4587), .B1(round_ctr_reg[0]), .Y(
        n3925) );
  INVX1 U1417 ( .A(n1732), .Y(n4587) );
  BUFX2 U1418 ( .A(n740), .Y(n4030) );
  BUFX2 U1419 ( .A(n740), .Y(n4031) );
  BUFX2 U1420 ( .A(n740), .Y(n4032) );
  BUFX2 U1421 ( .A(n740), .Y(n4033) );
  BUFX2 U1422 ( .A(n737), .Y(n4115) );
  BUFX2 U1423 ( .A(n736), .Y(n4143) );
  BUFX2 U1424 ( .A(n737), .Y(n4116) );
  BUFX2 U1425 ( .A(n736), .Y(n4144) );
  BUFX2 U1426 ( .A(n737), .Y(n4117) );
  BUFX2 U1427 ( .A(n736), .Y(n4145) );
  BUFX2 U1428 ( .A(n738), .Y(n4086) );
  BUFX2 U1429 ( .A(n739), .Y(n4059) );
  BUFX2 U1430 ( .A(n738), .Y(n4087) );
  BUFX2 U1431 ( .A(n739), .Y(n4060) );
  BUFX2 U1432 ( .A(n738), .Y(n4088) );
  BUFX2 U1433 ( .A(n739), .Y(n4061) );
  BUFX2 U1434 ( .A(n738), .Y(n4089) );
  BUFX2 U1435 ( .A(n729), .Y(n4283) );
  BUFX2 U1436 ( .A(n727), .Y(n4311) );
  BUFX2 U1437 ( .A(n729), .Y(n4284) );
  BUFX2 U1438 ( .A(n727), .Y(n4312) );
  BUFX2 U1439 ( .A(n729), .Y(n4285) );
  BUFX2 U1440 ( .A(n727), .Y(n4313) );
  BUFX2 U1441 ( .A(n735), .Y(n4171) );
  BUFX2 U1442 ( .A(n733), .Y(n4199) );
  BUFX2 U1443 ( .A(n735), .Y(n4172) );
  BUFX2 U1444 ( .A(n733), .Y(n4200) );
  BUFX2 U1445 ( .A(n735), .Y(n4173) );
  BUFX2 U1446 ( .A(n733), .Y(n4201) );
  XOR2X1 U1447 ( .A(n5220), .B(prev_key1_reg[115]), .Y(n5233) );
  XOR3X1 U1448 ( .A(prev_key1_reg[51]), .B(prev_key1_reg[83]), .C(n5233), .Y(
        n5244) );
  AOI222XL U1449 ( .A0(n1705), .A1(n827), .B0(key[107]), .B1(n1680), .C0(n1693), .C1(n828), .Y(n826) );
  INVX1 U1450 ( .A(n4961), .Y(n828) );
  INVX1 U1451 ( .A(n5247), .Y(n1177) );
  INVX1 U1452 ( .A(n5235), .Y(n1049) );
  INVX1 U1453 ( .A(n5227), .Y(n921) );
  AOI222XL U1454 ( .A0(n5759), .A1(n56), .B0(key[11]), .B1(n1688), .C0(n1699), 
        .C1(n5721), .Y(n1210) );
  INVX1 U1455 ( .A(n4984), .Y(n1209) );
  AOI222XL U1456 ( .A0(n1711), .A1(n1083), .B0(key[43]), .B1(n1684), .C0(n1698), .C1(n5722), .Y(n1082) );
  INVX1 U1457 ( .A(n4972), .Y(n1081) );
  AOI222XL U1458 ( .A0(n1708), .A1(n43), .B0(key[75]), .B1(n1690), .C0(n1695), 
        .C1(n5723), .Y(n954) );
  INVX1 U1459 ( .A(n4964), .Y(n953) );
  AO22X1 U1460 ( .A0(sboxw[11]), .A1(n1620), .B0(n1607), .B1(n4984), .Y(n4985)
         );
  AO22X1 U1461 ( .A0(prev_key1_reg[43]), .A1(n1619), .B0(n5668), .B1(n4972), 
        .Y(n4973) );
  AO22X1 U1462 ( .A0(prev_key1_reg[75]), .A1(n1618), .B0(n1603), .B1(n4964), 
        .Y(n4965) );
  AO22X1 U1463 ( .A0(n3965), .A1(n1444), .B0(\key_mem[1][19] ), .B1(n3983), 
        .Y(n1974) );
  AO22X1 U1464 ( .A0(n3969), .A1(n1476), .B0(\key_mem[1][51] ), .B1(n3987), 
        .Y(n1942) );
  AO22X1 U1465 ( .A0(n3972), .A1(n1508), .B0(\key_mem[1][83] ), .B1(n3988), 
        .Y(n1910) );
  AO22X1 U1466 ( .A0(n4035), .A1(n1444), .B0(\key_mem[13][19] ), .B1(n4050), 
        .Y(n3510) );
  AO22X1 U1467 ( .A0(n4091), .A1(n701), .B0(\key_mem[11][19] ), .B1(n4109), 
        .Y(n3254) );
  AO22X1 U1468 ( .A0(n4147), .A1(n701), .B0(\key_mem[9][19] ), .B1(n4171), .Y(
        n2998) );
  AO22X1 U1469 ( .A0(n4204), .A1(n701), .B0(\key_mem[7][19] ), .B1(n4221), .Y(
        n2742) );
  AO22X1 U1470 ( .A0(n4259), .A1(n701), .B0(\key_mem[5][19] ), .B1(n4284), .Y(
        n2486) );
  AO22X1 U1471 ( .A0(n4315), .A1(n701), .B0(\key_mem[3][19] ), .B1(n4333), .Y(
        n2230) );
  AO22X1 U1472 ( .A0(n4039), .A1(n1476), .B0(\key_mem[13][51] ), .B1(n4056), 
        .Y(n3478) );
  AO22X1 U1473 ( .A0(n4095), .A1(n669), .B0(\key_mem[11][51] ), .B1(n4107), 
        .Y(n3222) );
  AO22X1 U1474 ( .A0(n4151), .A1(n669), .B0(\key_mem[9][51] ), .B1(n4173), .Y(
        n2966) );
  AO22X1 U1475 ( .A0(n4207), .A1(n669), .B0(\key_mem[7][51] ), .B1(n4219), .Y(
        n2710) );
  AO22X1 U1476 ( .A0(n4263), .A1(n669), .B0(\key_mem[5][51] ), .B1(n4276), .Y(
        n2454) );
  AO22X1 U1477 ( .A0(n4319), .A1(n669), .B0(\key_mem[3][51] ), .B1(n4327), .Y(
        n2198) );
  AO22X1 U1478 ( .A0(n4042), .A1(n1508), .B0(\key_mem[13][83] ), .B1(n4051), 
        .Y(n3446) );
  AO22X1 U1479 ( .A0(n4098), .A1(n637), .B0(\key_mem[11][83] ), .B1(n4111), 
        .Y(n3190) );
  AO22X1 U1480 ( .A0(n4154), .A1(n637), .B0(\key_mem[9][83] ), .B1(n4170), .Y(
        n2934) );
  AO22X1 U1481 ( .A0(n4210), .A1(n637), .B0(\key_mem[7][83] ), .B1(n4226), .Y(
        n2678) );
  AO22X1 U1482 ( .A0(n4266), .A1(n637), .B0(\key_mem[5][83] ), .B1(n4282), .Y(
        n2422) );
  AO22X1 U1483 ( .A0(n4322), .A1(n637), .B0(\key_mem[3][83] ), .B1(n4329), .Y(
        n2166) );
  AO22X1 U1484 ( .A0(n3965), .A1(n1436), .B0(\key_mem[1][11] ), .B1(n3990), 
        .Y(n1982) );
  AO22X1 U1485 ( .A0(n3968), .A1(n1468), .B0(\key_mem[1][43] ), .B1(n3990), 
        .Y(n1950) );
  AO22X1 U1486 ( .A0(n3971), .A1(n1500), .B0(\key_mem[1][75] ), .B1(n3982), 
        .Y(n1918) );
  AO22X1 U1487 ( .A0(n3974), .A1(n1532), .B0(\key_mem[1][107] ), .B1(n3985), 
        .Y(n1886) );
  AO22X1 U1488 ( .A0(n4035), .A1(n1436), .B0(\key_mem[13][11] ), .B1(n4053), 
        .Y(n3518) );
  AO22X1 U1489 ( .A0(n4091), .A1(n709), .B0(\key_mem[11][11] ), .B1(n4113), 
        .Y(n3262) );
  AO22X1 U1490 ( .A0(n4147), .A1(n709), .B0(\key_mem[9][11] ), .B1(n4169), .Y(
        n3006) );
  AO22X1 U1491 ( .A0(n4204), .A1(n709), .B0(\key_mem[7][11] ), .B1(n4219), .Y(
        n2750) );
  AO22X1 U1492 ( .A0(n4259), .A1(n709), .B0(\key_mem[5][11] ), .B1(n4281), .Y(
        n2494) );
  AO22X1 U1493 ( .A0(n4315), .A1(n709), .B0(\key_mem[3][11] ), .B1(n4334), .Y(
        n2238) );
  AO22X1 U1494 ( .A0(n4038), .A1(n1468), .B0(\key_mem[13][43] ), .B1(n4055), 
        .Y(n3486) );
  AO22X1 U1495 ( .A0(n4094), .A1(n677), .B0(\key_mem[11][43] ), .B1(n4113), 
        .Y(n3230) );
  AO22X1 U1496 ( .A0(n4150), .A1(n677), .B0(\key_mem[9][43] ), .B1(n4162), .Y(
        n2974) );
  AO22X1 U1497 ( .A0(n4202), .A1(n677), .B0(\key_mem[7][43] ), .B1(n4218), .Y(
        n2718) );
  AO22X1 U1498 ( .A0(n4262), .A1(n677), .B0(\key_mem[5][43] ), .B1(n4283), .Y(
        n2462) );
  AO22X1 U1499 ( .A0(n4318), .A1(n677), .B0(\key_mem[3][43] ), .B1(n4330), .Y(
        n2206) );
  AO22X1 U1500 ( .A0(n4041), .A1(n1500), .B0(\key_mem[13][75] ), .B1(n4055), 
        .Y(n3454) );
  AO22X1 U1501 ( .A0(n4097), .A1(n645), .B0(\key_mem[11][75] ), .B1(n4112), 
        .Y(n3198) );
  AO22X1 U1502 ( .A0(n4153), .A1(n645), .B0(\key_mem[9][75] ), .B1(n4166), .Y(
        n2942) );
  AO22X1 U1503 ( .A0(n4209), .A1(n645), .B0(\key_mem[7][75] ), .B1(n4216), .Y(
        n2686) );
  AO22X1 U1504 ( .A0(n4265), .A1(n645), .B0(\key_mem[5][75] ), .B1(n4271), .Y(
        n2430) );
  AO22X1 U1505 ( .A0(n4321), .A1(n645), .B0(\key_mem[3][75] ), .B1(n4332), .Y(
        n2174) );
  AO22X1 U1506 ( .A0(n4044), .A1(n1532), .B0(\key_mem[13][107] ), .B1(n4058), 
        .Y(n3422) );
  AO22X1 U1507 ( .A0(n4100), .A1(n613), .B0(\key_mem[11][107] ), .B1(n4109), 
        .Y(n3166) );
  AO22X1 U1508 ( .A0(n4156), .A1(n613), .B0(\key_mem[9][107] ), .B1(n4160), 
        .Y(n2910) );
  AO22X1 U1509 ( .A0(n4212), .A1(n613), .B0(\key_mem[7][107] ), .B1(n4224), 
        .Y(n2654) );
  AO22X1 U1510 ( .A0(n4268), .A1(n613), .B0(\key_mem[5][107] ), .B1(n4271), 
        .Y(n2398) );
  AO22X1 U1511 ( .A0(n4324), .A1(n613), .B0(\key_mem[3][107] ), .B1(n4336), 
        .Y(n2142) );
  AO22X1 U1512 ( .A0(n4007), .A1(n1444), .B0(\key_mem[14][19] ), .B1(n4031), 
        .Y(n3638) );
  AO22X1 U1513 ( .A0(n4063), .A1(n1444), .B0(\key_mem[12][19] ), .B1(n4076), 
        .Y(n3382) );
  AO22X1 U1514 ( .A0(n4119), .A1(n1444), .B0(\key_mem[10][19] ), .B1(n4143), 
        .Y(n3126) );
  AO22X1 U1515 ( .A0(n4175), .A1(n1444), .B0(\key_mem[8][19] ), .B1(n4199), 
        .Y(n2870) );
  AO22X1 U1516 ( .A0(n4232), .A1(n1444), .B0(\key_mem[6][19] ), .B1(n4252), 
        .Y(n2614) );
  AO22X1 U1517 ( .A0(n4287), .A1(n1444), .B0(\key_mem[4][19] ), .B1(n4301), 
        .Y(n2358) );
  AO22X1 U1518 ( .A0(n4343), .A1(n1444), .B0(\key_mem[2][19] ), .B1(n4364), 
        .Y(n2102) );
  AO22X1 U1519 ( .A0(n3958), .A1(n1444), .B0(\key_mem[0][19] ), .B1(n1720), 
        .Y(n1846) );
  AO22X1 U1520 ( .A0(n4011), .A1(n1476), .B0(\key_mem[14][51] ), .B1(n4030), 
        .Y(n3606) );
  AO22X1 U1521 ( .A0(n4067), .A1(n1476), .B0(\key_mem[12][51] ), .B1(n4083), 
        .Y(n3350) );
  AO22X1 U1522 ( .A0(n4123), .A1(n1476), .B0(\key_mem[10][51] ), .B1(n4145), 
        .Y(n3094) );
  AO22X1 U1523 ( .A0(n4179), .A1(n1476), .B0(\key_mem[8][51] ), .B1(n4201), 
        .Y(n2838) );
  AO22X1 U1524 ( .A0(n4236), .A1(n1476), .B0(\key_mem[6][51] ), .B1(n4244), 
        .Y(n2582) );
  AO22X1 U1525 ( .A0(n4291), .A1(n1476), .B0(\key_mem[4][51] ), .B1(n4313), 
        .Y(n2326) );
  AO22X1 U1526 ( .A0(n4347), .A1(n1476), .B0(\key_mem[2][51] ), .B1(n4360), 
        .Y(n2070) );
  AO22X1 U1527 ( .A0(n3955), .A1(n1476), .B0(\key_mem[0][51] ), .B1(n3929), 
        .Y(n1814) );
  AO22X1 U1528 ( .A0(n4014), .A1(n1508), .B0(\key_mem[14][83] ), .B1(n4021), 
        .Y(n3574) );
  AO22X1 U1529 ( .A0(n4070), .A1(n1508), .B0(\key_mem[12][83] ), .B1(n4082), 
        .Y(n3318) );
  AO22X1 U1530 ( .A0(n4126), .A1(n1508), .B0(\key_mem[10][83] ), .B1(n4141), 
        .Y(n3062) );
  AO22X1 U1531 ( .A0(n4182), .A1(n1508), .B0(\key_mem[8][83] ), .B1(n4197), 
        .Y(n2806) );
  AO22X1 U1532 ( .A0(n4239), .A1(n1508), .B0(\key_mem[6][83] ), .B1(n4250), 
        .Y(n2550) );
  AO22X1 U1533 ( .A0(n4294), .A1(n1508), .B0(\key_mem[4][83] ), .B1(n4310), 
        .Y(n2294) );
  AO22X1 U1534 ( .A0(n4350), .A1(n1508), .B0(\key_mem[2][83] ), .B1(n4369), 
        .Y(n2038) );
  AO22X1 U1535 ( .A0(n3951), .A1(n1508), .B0(\key_mem[0][83] ), .B1(n3947), 
        .Y(n1782) );
  AO22X1 U1536 ( .A0(n4007), .A1(n1436), .B0(\key_mem[14][11] ), .B1(n4028), 
        .Y(n3646) );
  AO22X1 U1537 ( .A0(n4063), .A1(n1436), .B0(\key_mem[12][11] ), .B1(n4078), 
        .Y(n3390) );
  AO22X1 U1538 ( .A0(n4119), .A1(n1436), .B0(\key_mem[10][11] ), .B1(n4141), 
        .Y(n3134) );
  AO22X1 U1539 ( .A0(n4175), .A1(n1436), .B0(\key_mem[8][11] ), .B1(n4197), 
        .Y(n2878) );
  AO22X1 U1540 ( .A0(n4232), .A1(n1436), .B0(\key_mem[6][11] ), .B1(n4253), 
        .Y(n2622) );
  AO22X1 U1541 ( .A0(n4287), .A1(n1436), .B0(\key_mem[4][11] ), .B1(n4309), 
        .Y(n2366) );
  AO22X1 U1542 ( .A0(n4343), .A1(n1436), .B0(\key_mem[2][11] ), .B1(n4365), 
        .Y(n2110) );
  AO22X1 U1543 ( .A0(n3959), .A1(n1436), .B0(\key_mem[0][11] ), .B1(n1720), 
        .Y(n1854) );
  AO22X1 U1544 ( .A0(n4010), .A1(n1468), .B0(\key_mem[14][43] ), .B1(n4020), 
        .Y(n3614) );
  AO22X1 U1545 ( .A0(n4066), .A1(n1468), .B0(\key_mem[12][43] ), .B1(n4083), 
        .Y(n3358) );
  AO22X1 U1546 ( .A0(n4122), .A1(n1468), .B0(\key_mem[10][43] ), .B1(n4137), 
        .Y(n3102) );
  AO22X1 U1547 ( .A0(n4178), .A1(n1468), .B0(\key_mem[8][43] ), .B1(n4193), 
        .Y(n2846) );
  AO22X1 U1548 ( .A0(n4235), .A1(n1468), .B0(\key_mem[6][43] ), .B1(n4257), 
        .Y(n2590) );
  AO22X1 U1549 ( .A0(n4290), .A1(n1468), .B0(\key_mem[4][43] ), .B1(n4310), 
        .Y(n2334) );
  AO22X1 U1550 ( .A0(n4346), .A1(n1468), .B0(\key_mem[2][43] ), .B1(n4356), 
        .Y(n2078) );
  AO22X1 U1551 ( .A0(n3955), .A1(n1468), .B0(\key_mem[0][43] ), .B1(n3928), 
        .Y(n1822) );
  AO22X1 U1552 ( .A0(n4013), .A1(n1500), .B0(\key_mem[14][75] ), .B1(n4019), 
        .Y(n3582) );
  AO22X1 U1553 ( .A0(n4069), .A1(n1500), .B0(\key_mem[12][75] ), .B1(n4075), 
        .Y(n3326) );
  AO22X1 U1554 ( .A0(n4125), .A1(n1500), .B0(\key_mem[10][75] ), .B1(n4134), 
        .Y(n3070) );
  AO22X1 U1555 ( .A0(n4181), .A1(n1500), .B0(\key_mem[8][75] ), .B1(n4191), 
        .Y(n2814) );
  AO22X1 U1556 ( .A0(n4238), .A1(n1500), .B0(\key_mem[6][75] ), .B1(n4251), 
        .Y(n2558) );
  AO22X1 U1557 ( .A0(n4293), .A1(n1500), .B0(\key_mem[4][75] ), .B1(n4310), 
        .Y(n2302) );
  AO22X1 U1558 ( .A0(n4349), .A1(n1500), .B0(\key_mem[2][75] ), .B1(n4366), 
        .Y(n2046) );
  AO22X1 U1559 ( .A0(n3952), .A1(n1500), .B0(\key_mem[0][75] ), .B1(n3931), 
        .Y(n1790) );
  AO22X1 U1560 ( .A0(n4016), .A1(n1532), .B0(\key_mem[14][107] ), .B1(n4029), 
        .Y(n3550) );
  AO22X1 U1561 ( .A0(n4072), .A1(n1532), .B0(\key_mem[12][107] ), .B1(n4084), 
        .Y(n3294) );
  AO22X1 U1562 ( .A0(n4128), .A1(n1532), .B0(\key_mem[10][107] ), .B1(n4131), 
        .Y(n3038) );
  AO22X1 U1563 ( .A0(n4184), .A1(n1532), .B0(\key_mem[8][107] ), .B1(n4187), 
        .Y(n2782) );
  AO22X1 U1564 ( .A0(n4241), .A1(n1532), .B0(\key_mem[6][107] ), .B1(n4250), 
        .Y(n2526) );
  AO22X1 U1565 ( .A0(n4296), .A1(n1532), .B0(\key_mem[4][107] ), .B1(n4309), 
        .Y(n2270) );
  AO22X1 U1566 ( .A0(n4352), .A1(n1532), .B0(\key_mem[2][107] ), .B1(n4359), 
        .Y(n2014) );
  AO22X1 U1567 ( .A0(n3949), .A1(n1532), .B0(\key_mem[0][107] ), .B1(n1717), 
        .Y(n1758) );
  XNOR2X1 U1568 ( .A(n5244), .B(sboxw[19]), .Y(n7) );
  OAI221XL U1569 ( .A0(n1668), .A1(n4962), .B0(n4961), .B1(n1657), .C0(n4960), 
        .Y(n3805) );
  INVX1 U1570 ( .A(key[107]), .Y(n4962) );
  AOI221XL U1571 ( .A0(n1642), .A1(n827), .B0(n1634), .B1(key[235]), .C0(n4959), .Y(n4960) );
  AO22X1 U1572 ( .A0(prev_key1_reg[107]), .A1(n1617), .B0(n1605), .B1(n4958), 
        .Y(n4959) );
  OAI221XL U1573 ( .A0(n1668), .A1(n4988), .B0(n1663), .B1(n4987), .C0(n4986), 
        .Y(n3901) );
  INVX1 U1574 ( .A(key[11]), .Y(n4988) );
  INVX1 U1575 ( .A(n5721), .Y(n4987) );
  AOI221XL U1576 ( .A0(n1642), .A1(n56), .B0(n1635), .B1(key[139]), .C0(n4985), 
        .Y(n4986) );
  OAI221XL U1577 ( .A0(n1669), .A1(n5251), .B0(n1651), .B1(n5250), .C0(n5249), 
        .Y(n3893) );
  INVX1 U1578 ( .A(key[19]), .Y(n5251) );
  AOI221XL U1579 ( .A0(n1638), .A1(n7), .B0(n1627), .B1(key[147]), .C0(n5248), 
        .Y(n5249) );
  OAI221XL U1580 ( .A0(n1668), .A1(n4976), .B0(n1662), .B1(n4975), .C0(n4974), 
        .Y(n3869) );
  INVX1 U1581 ( .A(key[43]), .Y(n4976) );
  INVX1 U1582 ( .A(n5722), .Y(n4975) );
  AOI221XL U1583 ( .A0(n1642), .A1(n1083), .B0(n1635), .B1(key[171]), .C0(
        n4973), .Y(n4974) );
  OAI221XL U1584 ( .A0(n1669), .A1(n5239), .B0(n1651), .B1(n5238), .C0(n5237), 
        .Y(n3861) );
  INVX1 U1585 ( .A(key[51]), .Y(n5239) );
  AOI221XL U1586 ( .A0(n1638), .A1(n1051), .B0(n1627), .B1(key[179]), .C0(
        n5236), .Y(n5237) );
  OAI221XL U1587 ( .A0(n1668), .A1(n4968), .B0(n1663), .B1(n4967), .C0(n4966), 
        .Y(n3837) );
  INVX1 U1588 ( .A(key[75]), .Y(n4968) );
  INVX1 U1589 ( .A(n5723), .Y(n4967) );
  AOI221XL U1590 ( .A0(n1642), .A1(n43), .B0(n1631), .B1(key[203]), .C0(n4965), 
        .Y(n4966) );
  OAI221XL U1591 ( .A0(n1669), .A1(n5231), .B0(n1651), .B1(n5230), .C0(n5229), 
        .Y(n3829) );
  INVX1 U1592 ( .A(key[83]), .Y(n5231) );
  AOI221XL U1593 ( .A0(n1639), .A1(n6), .B0(n1627), .B1(key[211]), .C0(n5228), 
        .Y(n5229) );
  XOR2X1 U1594 ( .A(n5056), .B(prev_key1_reg[110]), .Y(n5068) );
  XOR2X1 U1595 ( .A(n4858), .B(prev_key1_reg[104]), .Y(n4871) );
  INVX1 U1596 ( .A(n5082), .Y(n1197) );
  XOR2X1 U1597 ( .A(n5056), .B(prev_key0_reg[110]), .Y(n5060) );
  OAI221XL U1598 ( .A0(n965), .A1(n3995), .B0(n3942), .B1(n5785), .C0(n966), 
        .Y(n648) );
  OAI221XL U1599 ( .A0(n1666), .A1(n4614), .B0(n1653), .B1(n4613), .C0(n4612), 
        .Y(n3848) );
  INVX1 U1600 ( .A(key[64]), .Y(n4614) );
  INVX1 U1601 ( .A(n5756), .Y(n4613) );
  AOI221XL U1602 ( .A0(n1647), .A1(n35), .B0(n1622), .B1(key[192]), .C0(n4611), 
        .Y(n4612) );
  XOR3X1 U1603 ( .A(prev_key1_reg[46]), .B(prev_key1_reg[78]), .C(n5068), .Y(
        n5079) );
  XOR3X1 U1604 ( .A(prev_key1_reg[40]), .B(prev_key1_reg[72]), .C(n4871), .Y(
        n4882) );
  AOI222XL U1605 ( .A0(n1706), .A1(n871), .B0(key[96]), .B1(n1681), .C0(n1694), 
        .C1(n872), .Y(n870) );
  INVX1 U1606 ( .A(n4607), .Y(n872) );
  AOI222XL U1607 ( .A0(n5759), .A1(n53), .B0(key[6]), .B1(n1688), .C0(n1701), 
        .C1(n5736), .Y(n1230) );
  INVX1 U1608 ( .A(n4820), .Y(n1229) );
  AOI222XL U1609 ( .A0(n1716), .A1(n1127), .B0(key[32]), .B1(n1686), .C0(n1701), .C1(n5755), .Y(n1126) );
  AOI222XL U1610 ( .A0(n1714), .A1(n1103), .B0(key[38]), .B1(n1684), .C0(n5758), .C1(n5737), .Y(n1102) );
  INVX1 U1611 ( .A(n4808), .Y(n1101) );
  AOI222XL U1612 ( .A0(n1709), .A1(n35), .B0(key[64]), .B1(n5757), .C0(n1696), 
        .C1(n5756), .Y(n998) );
  AOI222XL U1613 ( .A0(n1708), .A1(n40), .B0(key[70]), .B1(n1685), .C0(n1695), 
        .C1(n5738), .Y(n974) );
  INVX1 U1614 ( .A(n4800), .Y(n973) );
  XNOR2X1 U1615 ( .A(n5068), .B(prev_key1_reg[78]), .Y(n8) );
  OAI221XL U1616 ( .A0(n1093), .A1(n4004), .B0(n3939), .B1(n5787), .C0(n1094), 
        .Y(n680) );
  OAI221XL U1617 ( .A0(n1069), .A1(n4004), .B0(n3939), .B1(n5867), .C0(n1070), 
        .Y(n674) );
  INVX1 U1618 ( .A(n5070), .Y(n1069) );
  AO22X1 U1619 ( .A0(sboxw[6]), .A1(n1617), .B0(n1606), .B1(n4820), .Y(n4821)
         );
  AO22X1 U1620 ( .A0(prev_key1_reg[38]), .A1(n1618), .B0(n1607), .B1(n4808), 
        .Y(n4809) );
  AO22X1 U1621 ( .A0(prev_key1_reg[70]), .A1(n1617), .B0(n1606), .B1(n4800), 
        .Y(n4801) );
  AOI222XL U1622 ( .A0(n1704), .A1(n815), .B0(key[110]), .B1(n1679), .C0(n1692), .C1(n816), .Y(n814) );
  INVX1 U1623 ( .A(n5060), .Y(n816) );
  AO22X1 U1624 ( .A0(n3964), .A1(n1431), .B0(\key_mem[1][6] ), .B1(n3991), .Y(
        n1987) );
  AO22X1 U1625 ( .A0(n3964), .A1(n1433), .B0(\key_mem[1][8] ), .B1(n3982), .Y(
        n1985) );
  AO22X1 U1626 ( .A0(n3965), .A1(n1439), .B0(\key_mem[1][14] ), .B1(n3983), 
        .Y(n1979) );
  AO22X1 U1627 ( .A0(n3967), .A1(n1457), .B0(\key_mem[1][32] ), .B1(n3990), 
        .Y(n1961) );
  AO22X1 U1628 ( .A0(n3967), .A1(n1463), .B0(\key_mem[1][38] ), .B1(n3991), 
        .Y(n1955) );
  AO22X1 U1629 ( .A0(n3970), .A1(n1489), .B0(\key_mem[1][64] ), .B1(n3987), 
        .Y(n1929) );
  AO22X1 U1630 ( .A0(n3971), .A1(n1495), .B0(\key_mem[1][70] ), .B1(n3981), 
        .Y(n1923) );
  AO22X1 U1631 ( .A0(n3973), .A1(n1521), .B0(\key_mem[1][96] ), .B1(n3985), 
        .Y(n1897) );
  AO22X1 U1632 ( .A0(n3975), .A1(n1535), .B0(\key_mem[1][110] ), .B1(n3988), 
        .Y(n1883) );
  AO22X1 U1633 ( .A0(n3975), .A1(n1540), .B0(\key_mem[1][115] ), .B1(n3987), 
        .Y(n1878) );
  AO22X1 U1634 ( .A0(n4034), .A1(n1431), .B0(\key_mem[13][6] ), .B1(n4052), 
        .Y(n3523) );
  AO22X1 U1635 ( .A0(n4090), .A1(n714), .B0(\key_mem[11][6] ), .B1(n4108), .Y(
        n3267) );
  AO22X1 U1636 ( .A0(n4146), .A1(n714), .B0(\key_mem[9][6] ), .B1(n4164), .Y(
        n3011) );
  AO22X1 U1637 ( .A0(n4203), .A1(n714), .B0(\key_mem[7][6] ), .B1(n4217), .Y(
        n2755) );
  AO22X1 U1638 ( .A0(n4258), .A1(n714), .B0(\key_mem[5][6] ), .B1(n4276), .Y(
        n2499) );
  AO22X1 U1639 ( .A0(n4314), .A1(n714), .B0(\key_mem[3][6] ), .B1(n4332), .Y(
        n2243) );
  AO22X1 U1640 ( .A0(n4034), .A1(n1433), .B0(\key_mem[13][8] ), .B1(n4054), 
        .Y(n3521) );
  AO22X1 U1641 ( .A0(n4090), .A1(n712), .B0(\key_mem[11][8] ), .B1(n4110), .Y(
        n3265) );
  AO22X1 U1642 ( .A0(n4146), .A1(n712), .B0(\key_mem[9][8] ), .B1(n4166), .Y(
        n3009) );
  AO22X1 U1643 ( .A0(n4203), .A1(n712), .B0(\key_mem[7][8] ), .B1(n4216), .Y(
        n2753) );
  AO22X1 U1644 ( .A0(n4258), .A1(n712), .B0(\key_mem[5][8] ), .B1(n4278), .Y(
        n2497) );
  AO22X1 U1645 ( .A0(n4314), .A1(n712), .B0(\key_mem[3][8] ), .B1(n4334), .Y(
        n2241) );
  AO22X1 U1646 ( .A0(n4035), .A1(n1439), .B0(\key_mem[13][14] ), .B1(n4047), 
        .Y(n3515) );
  AO22X1 U1647 ( .A0(n4091), .A1(n706), .B0(\key_mem[11][14] ), .B1(n4106), 
        .Y(n3259) );
  AO22X1 U1648 ( .A0(n4147), .A1(n706), .B0(\key_mem[9][14] ), .B1(n4160), .Y(
        n3003) );
  AO22X1 U1649 ( .A0(n4204), .A1(n706), .B0(\key_mem[7][14] ), .B1(n4221), .Y(
        n2747) );
  AO22X1 U1650 ( .A0(n4259), .A1(n706), .B0(\key_mem[5][14] ), .B1(n4279), .Y(
        n2491) );
  AO22X1 U1651 ( .A0(n4315), .A1(n706), .B0(\key_mem[3][14] ), .B1(n4337), .Y(
        n2235) );
  AO22X1 U1652 ( .A0(n4037), .A1(n1457), .B0(\key_mem[13][32] ), .B1(n4054), 
        .Y(n3497) );
  AO22X1 U1653 ( .A0(n4093), .A1(n688), .B0(\key_mem[11][32] ), .B1(n4105), 
        .Y(n3241) );
  AO22X1 U1654 ( .A0(n4149), .A1(n688), .B0(\key_mem[9][32] ), .B1(n4172), .Y(
        n2985) );
  AO22X1 U1655 ( .A0(n4206), .A1(n688), .B0(\key_mem[7][32] ), .B1(n4222), .Y(
        n2729) );
  AO22X1 U1656 ( .A0(n4261), .A1(n688), .B0(\key_mem[5][32] ), .B1(n4284), .Y(
        n2473) );
  AO22X1 U1657 ( .A0(n4317), .A1(n688), .B0(\key_mem[3][32] ), .B1(n4335), .Y(
        n2217) );
  AO22X1 U1658 ( .A0(n4037), .A1(n1463), .B0(\key_mem[13][38] ), .B1(n4047), 
        .Y(n3491) );
  AO22X1 U1659 ( .A0(n4093), .A1(n682), .B0(\key_mem[11][38] ), .B1(n4117), 
        .Y(n3235) );
  AO22X1 U1660 ( .A0(n4149), .A1(n682), .B0(\key_mem[9][38] ), .B1(n4171), .Y(
        n2979) );
  AO22X1 U1661 ( .A0(n4206), .A1(n682), .B0(\key_mem[7][38] ), .B1(n4223), .Y(
        n2723) );
  AO22X1 U1662 ( .A0(n4261), .A1(n682), .B0(\key_mem[5][38] ), .B1(n4275), .Y(
        n2467) );
  AO22X1 U1663 ( .A0(n4317), .A1(n682), .B0(\key_mem[3][38] ), .B1(n4334), .Y(
        n2211) );
  AO22X1 U1664 ( .A0(n4040), .A1(n1489), .B0(\key_mem[13][64] ), .B1(n4056), 
        .Y(n3465) );
  AO22X1 U1665 ( .A0(n4096), .A1(n656), .B0(\key_mem[11][64] ), .B1(n4114), 
        .Y(n3209) );
  AO22X1 U1666 ( .A0(n4152), .A1(n656), .B0(\key_mem[9][64] ), .B1(n4163), .Y(
        n2953) );
  AO22X1 U1667 ( .A0(n4208), .A1(n656), .B0(\key_mem[7][64] ), .B1(n4219), .Y(
        n2697) );
  AO22X1 U1668 ( .A0(n4264), .A1(n656), .B0(\key_mem[5][64] ), .B1(n4276), .Y(
        n2441) );
  AO22X1 U1669 ( .A0(n4320), .A1(n656), .B0(\key_mem[3][64] ), .B1(n4327), .Y(
        n2185) );
  AO22X1 U1670 ( .A0(n4041), .A1(n1495), .B0(\key_mem[13][70] ), .B1(n4050), 
        .Y(n3459) );
  AO22X1 U1671 ( .A0(n4097), .A1(n650), .B0(\key_mem[11][70] ), .B1(n4114), 
        .Y(n3203) );
  AO22X1 U1672 ( .A0(n4153), .A1(n650), .B0(\key_mem[9][70] ), .B1(n4162), .Y(
        n2947) );
  AO22X1 U1673 ( .A0(n4209), .A1(n650), .B0(\key_mem[7][70] ), .B1(n4214), .Y(
        n2691) );
  AO22X1 U1674 ( .A0(n4265), .A1(n650), .B0(\key_mem[5][70] ), .B1(n4275), .Y(
        n2435) );
  AO22X1 U1675 ( .A0(n4321), .A1(n650), .B0(\key_mem[3][70] ), .B1(n4328), .Y(
        n2179) );
  AO22X1 U1676 ( .A0(n4043), .A1(n1521), .B0(\key_mem[13][96] ), .B1(n4057), 
        .Y(n3433) );
  AO22X1 U1677 ( .A0(n4099), .A1(n624), .B0(\key_mem[11][96] ), .B1(n4109), 
        .Y(n3177) );
  AO22X1 U1678 ( .A0(n4155), .A1(n624), .B0(\key_mem[9][96] ), .B1(n4168), .Y(
        n2921) );
  AO22X1 U1679 ( .A0(n4211), .A1(n624), .B0(\key_mem[7][96] ), .B1(n4216), .Y(
        n2665) );
  AO22X1 U1680 ( .A0(n4267), .A1(n624), .B0(\key_mem[5][96] ), .B1(n4280), .Y(
        n2409) );
  AO22X1 U1681 ( .A0(n4323), .A1(n624), .B0(\key_mem[3][96] ), .B1(n4335), .Y(
        n2153) );
  AO22X1 U1682 ( .A0(n4045), .A1(n1535), .B0(\key_mem[13][110] ), .B1(n4052), 
        .Y(n3419) );
  AO22X1 U1683 ( .A0(n4101), .A1(n610), .B0(\key_mem[11][110] ), .B1(n4103), 
        .Y(n3163) );
  AO22X1 U1684 ( .A0(n4157), .A1(n610), .B0(\key_mem[9][110] ), .B1(n4170), 
        .Y(n2907) );
  AO22X1 U1685 ( .A0(n4213), .A1(n610), .B0(\key_mem[7][110] ), .B1(n4224), 
        .Y(n2651) );
  AO22X1 U1686 ( .A0(n4269), .A1(n610), .B0(\key_mem[5][110] ), .B1(n4282), 
        .Y(n2395) );
  AO22X1 U1687 ( .A0(n4325), .A1(n610), .B0(\key_mem[3][110] ), .B1(n4336), 
        .Y(n2139) );
  AO22X1 U1688 ( .A0(n4045), .A1(n1540), .B0(\key_mem[13][115] ), .B1(n4058), 
        .Y(n3414) );
  AO22X1 U1689 ( .A0(n4101), .A1(n605), .B0(\key_mem[11][115] ), .B1(n4112), 
        .Y(n3158) );
  AO22X1 U1690 ( .A0(n4157), .A1(n605), .B0(\key_mem[9][115] ), .B1(n4161), 
        .Y(n2902) );
  AO22X1 U1691 ( .A0(n4213), .A1(n605), .B0(\key_mem[7][115] ), .B1(n4225), 
        .Y(n2646) );
  AO22X1 U1692 ( .A0(n4269), .A1(n605), .B0(\key_mem[5][115] ), .B1(n4272), 
        .Y(n2390) );
  AO22X1 U1693 ( .A0(n4325), .A1(n605), .B0(\key_mem[3][115] ), .B1(n4338), 
        .Y(n2134) );
  AO22X1 U1694 ( .A0(n4006), .A1(n1431), .B0(\key_mem[14][6] ), .B1(n4024), 
        .Y(n3651) );
  AO22X1 U1695 ( .A0(n4062), .A1(n1431), .B0(\key_mem[12][6] ), .B1(n4080), 
        .Y(n3395) );
  AO22X1 U1696 ( .A0(n4118), .A1(n1431), .B0(\key_mem[10][6] ), .B1(n4136), 
        .Y(n3139) );
  AO22X1 U1697 ( .A0(n4174), .A1(n1431), .B0(\key_mem[8][6] ), .B1(n4192), .Y(
        n2883) );
  AO22X1 U1698 ( .A0(n4231), .A1(n1431), .B0(\key_mem[6][6] ), .B1(n4250), .Y(
        n2627) );
  AO22X1 U1699 ( .A0(n4286), .A1(n1431), .B0(\key_mem[4][6] ), .B1(n4304), .Y(
        n2371) );
  AO22X1 U1700 ( .A0(n4342), .A1(n1431), .B0(\key_mem[2][6] ), .B1(n4360), .Y(
        n2115) );
  AO22X1 U1701 ( .A0(n3959), .A1(n1431), .B0(\key_mem[0][6] ), .B1(n1719), .Y(
        n1859) );
  AO22X1 U1702 ( .A0(n4006), .A1(n1433), .B0(\key_mem[14][8] ), .B1(n4025), 
        .Y(n3649) );
  AO22X1 U1703 ( .A0(n4062), .A1(n1433), .B0(\key_mem[12][8] ), .B1(n4082), 
        .Y(n3393) );
  AO22X1 U1704 ( .A0(n4118), .A1(n1433), .B0(\key_mem[10][8] ), .B1(n4138), 
        .Y(n3137) );
  AO22X1 U1705 ( .A0(n4174), .A1(n1433), .B0(\key_mem[8][8] ), .B1(n4194), .Y(
        n2881) );
  AO22X1 U1706 ( .A0(n4231), .A1(n1433), .B0(\key_mem[6][8] ), .B1(n4252), .Y(
        n2625) );
  AO22X1 U1707 ( .A0(n4286), .A1(n1433), .B0(\key_mem[4][8] ), .B1(n4306), .Y(
        n2369) );
  AO22X1 U1708 ( .A0(n4342), .A1(n1433), .B0(\key_mem[2][8] ), .B1(n4362), .Y(
        n2113) );
  AO22X1 U1709 ( .A0(n3959), .A1(n1433), .B0(\key_mem[0][8] ), .B1(n1719), .Y(
        n1857) );
  AO22X1 U1710 ( .A0(n4007), .A1(n1439), .B0(\key_mem[14][14] ), .B1(n4024), 
        .Y(n3643) );
  AO22X1 U1711 ( .A0(n4063), .A1(n1439), .B0(\key_mem[12][14] ), .B1(n4080), 
        .Y(n3387) );
  AO22X1 U1712 ( .A0(n4119), .A1(n1439), .B0(\key_mem[10][14] ), .B1(n4131), 
        .Y(n3131) );
  AO22X1 U1713 ( .A0(n4175), .A1(n1439), .B0(\key_mem[8][14] ), .B1(n4187), 
        .Y(n2875) );
  AO22X1 U1714 ( .A0(n4232), .A1(n1439), .B0(\key_mem[6][14] ), .B1(n4254), 
        .Y(n2619) );
  AO22X1 U1715 ( .A0(n4287), .A1(n1439), .B0(\key_mem[4][14] ), .B1(n4312), 
        .Y(n2363) );
  AO22X1 U1716 ( .A0(n4343), .A1(n1439), .B0(\key_mem[2][14] ), .B1(n4358), 
        .Y(n2107) );
  AO22X1 U1717 ( .A0(n3958), .A1(n1439), .B0(\key_mem[0][14] ), .B1(n1720), 
        .Y(n1851) );
  AO22X1 U1718 ( .A0(n4009), .A1(n1457), .B0(\key_mem[14][32] ), .B1(n4033), 
        .Y(n3625) );
  AO22X1 U1719 ( .A0(n4065), .A1(n1457), .B0(\key_mem[12][32] ), .B1(n4088), 
        .Y(n3369) );
  AO22X1 U1720 ( .A0(n4121), .A1(n1457), .B0(\key_mem[10][32] ), .B1(n4144), 
        .Y(n3113) );
  AO22X1 U1721 ( .A0(n4177), .A1(n1457), .B0(\key_mem[8][32] ), .B1(n4200), 
        .Y(n2857) );
  AO22X1 U1722 ( .A0(n4234), .A1(n1457), .B0(\key_mem[6][32] ), .B1(n4255), 
        .Y(n2601) );
  AO22X1 U1723 ( .A0(n4289), .A1(n1457), .B0(\key_mem[4][32] ), .B1(n4300), 
        .Y(n2345) );
  AO22X1 U1724 ( .A0(n4345), .A1(n1457), .B0(\key_mem[2][32] ), .B1(n4363), 
        .Y(n2089) );
  AO22X1 U1725 ( .A0(n3957), .A1(n1457), .B0(\key_mem[0][32] ), .B1(n1736), 
        .Y(n1833) );
  AO22X1 U1726 ( .A0(n4009), .A1(n1463), .B0(\key_mem[14][38] ), .B1(n4027), 
        .Y(n3619) );
  AO22X1 U1727 ( .A0(n4065), .A1(n1463), .B0(\key_mem[12][38] ), .B1(n4086), 
        .Y(n3363) );
  AO22X1 U1728 ( .A0(n4121), .A1(n1463), .B0(\key_mem[10][38] ), .B1(n4143), 
        .Y(n3107) );
  AO22X1 U1729 ( .A0(n4177), .A1(n1463), .B0(\key_mem[8][38] ), .B1(n4199), 
        .Y(n2851) );
  AO22X1 U1730 ( .A0(n4234), .A1(n1463), .B0(\key_mem[6][38] ), .B1(n4256), 
        .Y(n2595) );
  AO22X1 U1731 ( .A0(n4289), .A1(n1463), .B0(\key_mem[4][38] ), .B1(n4301), 
        .Y(n2339) );
  AO22X1 U1732 ( .A0(n4345), .A1(n1463), .B0(\key_mem[2][38] ), .B1(n4362), 
        .Y(n2083) );
  AO22X1 U1733 ( .A0(n3956), .A1(n1463), .B0(\key_mem[0][38] ), .B1(n1736), 
        .Y(n1827) );
  AO22X1 U1734 ( .A0(n4012), .A1(n1489), .B0(\key_mem[14][64] ), .B1(n4031), 
        .Y(n3593) );
  AO22X1 U1735 ( .A0(n4068), .A1(n1489), .B0(\key_mem[12][64] ), .B1(n4080), 
        .Y(n3337) );
  AO22X1 U1736 ( .A0(n4124), .A1(n1489), .B0(\key_mem[10][64] ), .B1(n4139), 
        .Y(n3081) );
  AO22X1 U1737 ( .A0(n4180), .A1(n1489), .B0(\key_mem[8][64] ), .B1(n4195), 
        .Y(n2825) );
  AO22X1 U1738 ( .A0(n4237), .A1(n1489), .B0(\key_mem[6][64] ), .B1(n4254), 
        .Y(n2569) );
  AO22X1 U1739 ( .A0(n4292), .A1(n1489), .B0(\key_mem[4][64] ), .B1(n4299), 
        .Y(n2313) );
  AO22X1 U1740 ( .A0(n4348), .A1(n1489), .B0(\key_mem[2][64] ), .B1(n4367), 
        .Y(n2057) );
  AO22X1 U1741 ( .A0(n3953), .A1(n1489), .B0(\key_mem[0][64] ), .B1(n3930), 
        .Y(n1801) );
  AO22X1 U1742 ( .A0(n4013), .A1(n1495), .B0(\key_mem[14][70] ), .B1(n4025), 
        .Y(n3587) );
  AO22X1 U1743 ( .A0(n4069), .A1(n1495), .B0(\key_mem[12][70] ), .B1(n4079), 
        .Y(n3331) );
  AO22X1 U1744 ( .A0(n4125), .A1(n1495), .B0(\key_mem[10][70] ), .B1(n4138), 
        .Y(n3075) );
  AO22X1 U1745 ( .A0(n4181), .A1(n1495), .B0(\key_mem[8][70] ), .B1(n4194), 
        .Y(n2819) );
  AO22X1 U1746 ( .A0(n4238), .A1(n1495), .B0(\key_mem[6][70] ), .B1(n4249), 
        .Y(n2563) );
  AO22X1 U1747 ( .A0(n4293), .A1(n1495), .B0(\key_mem[4][70] ), .B1(n4310), 
        .Y(n2307) );
  AO22X1 U1748 ( .A0(n4349), .A1(n1495), .B0(\key_mem[2][70] ), .B1(n4368), 
        .Y(n2051) );
  AO22X1 U1749 ( .A0(n3953), .A1(n1495), .B0(\key_mem[0][70] ), .B1(n3931), 
        .Y(n1795) );
  AO22X1 U1750 ( .A0(n4015), .A1(n1521), .B0(\key_mem[14][96] ), .B1(n4026), 
        .Y(n3561) );
  AO22X1 U1751 ( .A0(n4071), .A1(n1521), .B0(\key_mem[12][96] ), .B1(n4079), 
        .Y(n3305) );
  AO22X1 U1752 ( .A0(n4127), .A1(n1521), .B0(\key_mem[10][96] ), .B1(n4142), 
        .Y(n3049) );
  AO22X1 U1753 ( .A0(n4183), .A1(n1521), .B0(\key_mem[8][96] ), .B1(n4198), 
        .Y(n2793) );
  AO22X1 U1754 ( .A0(n4240), .A1(n1521), .B0(\key_mem[6][96] ), .B1(n4245), 
        .Y(n2537) );
  AO22X1 U1755 ( .A0(n4295), .A1(n1521), .B0(\key_mem[4][96] ), .B1(n4310), 
        .Y(n2281) );
  AO22X1 U1756 ( .A0(n4351), .A1(n1521), .B0(\key_mem[2][96] ), .B1(n4364), 
        .Y(n2025) );
  AO22X1 U1757 ( .A0(n3950), .A1(n1521), .B0(\key_mem[0][96] ), .B1(n3932), 
        .Y(n1769) );
  AO22X1 U1758 ( .A0(n4017), .A1(n1535), .B0(\key_mem[14][110] ), .B1(n4028), 
        .Y(n3547) );
  AO22X1 U1759 ( .A0(n4073), .A1(n1535), .B0(\key_mem[12][110] ), .B1(n4084), 
        .Y(n3291) );
  AO22X1 U1760 ( .A0(n4129), .A1(n1535), .B0(\key_mem[10][110] ), .B1(n4142), 
        .Y(n3035) );
  AO22X1 U1761 ( .A0(n4185), .A1(n1535), .B0(\key_mem[8][110] ), .B1(n4198), 
        .Y(n2779) );
  AO22X1 U1762 ( .A0(n4242), .A1(n1535), .B0(\key_mem[6][110] ), .B1(n4249), 
        .Y(n2523) );
  AO22X1 U1763 ( .A0(n4297), .A1(n1535), .B0(\key_mem[4][110] ), .B1(n4308), 
        .Y(n2267) );
  AO22X1 U1764 ( .A0(n4353), .A1(n1535), .B0(\key_mem[2][110] ), .B1(n4357), 
        .Y(n2011) );
  AO22X1 U1765 ( .A0(n3949), .A1(n1535), .B0(\key_mem[0][110] ), .B1(n3933), 
        .Y(n1755) );
  AO22X1 U1766 ( .A0(n4017), .A1(n1540), .B0(\key_mem[14][115] ), .B1(n740), 
        .Y(n3542) );
  AO22X1 U1767 ( .A0(n4073), .A1(n1540), .B0(\key_mem[12][115] ), .B1(n4085), 
        .Y(n3286) );
  AO22X1 U1768 ( .A0(n4129), .A1(n1540), .B0(\key_mem[10][115] ), .B1(n4132), 
        .Y(n3030) );
  AO22X1 U1769 ( .A0(n4185), .A1(n1540), .B0(\key_mem[8][115] ), .B1(n4188), 
        .Y(n2774) );
  AO22X1 U1770 ( .A0(n4242), .A1(n1540), .B0(\key_mem[6][115] ), .B1(n4253), 
        .Y(n2518) );
  AO22X1 U1771 ( .A0(n4297), .A1(n1540), .B0(\key_mem[4][115] ), .B1(n4309), 
        .Y(n2262) );
  AO22X1 U1772 ( .A0(n4353), .A1(n1540), .B0(\key_mem[2][115] ), .B1(n4358), 
        .Y(n2006) );
  AO22X1 U1773 ( .A0(n3948), .A1(n1540), .B0(\key_mem[0][115] ), .B1(n3933), 
        .Y(n1750) );
  AO22X1 U1774 ( .A0(n3968), .A1(n1465), .B0(\key_mem[1][40] ), .B1(n3987), 
        .Y(n1953) );
  AO22X1 U1775 ( .A0(n3968), .A1(n1471), .B0(\key_mem[1][46] ), .B1(n3985), 
        .Y(n1947) );
  AO22X1 U1776 ( .A0(n4038), .A1(n1465), .B0(\key_mem[13][40] ), .B1(n4059), 
        .Y(n3489) );
  AO22X1 U1777 ( .A0(n4094), .A1(n680), .B0(\key_mem[11][40] ), .B1(n4110), 
        .Y(n3233) );
  AO22X1 U1778 ( .A0(n4150), .A1(n680), .B0(\key_mem[9][40] ), .B1(n4164), .Y(
        n2977) );
  AO22X1 U1779 ( .A0(n4202), .A1(n680), .B0(\key_mem[7][40] ), .B1(n4223), .Y(
        n2721) );
  AO22X1 U1780 ( .A0(n4262), .A1(n680), .B0(\key_mem[5][40] ), .B1(n4275), .Y(
        n2465) );
  AO22X1 U1781 ( .A0(n4318), .A1(n680), .B0(\key_mem[3][40] ), .B1(n4330), .Y(
        n2209) );
  AO22X1 U1782 ( .A0(n4038), .A1(n1471), .B0(\key_mem[13][46] ), .B1(n4047), 
        .Y(n3483) );
  AO22X1 U1783 ( .A0(n4094), .A1(n674), .B0(\key_mem[11][46] ), .B1(n4111), 
        .Y(n3227) );
  AO22X1 U1784 ( .A0(n4150), .A1(n674), .B0(\key_mem[9][46] ), .B1(n4159), .Y(
        n2971) );
  AO22X1 U1785 ( .A0(n732), .A1(n674), .B0(\key_mem[7][46] ), .B1(n4214), .Y(
        n2715) );
  AO22X1 U1786 ( .A0(n4262), .A1(n674), .B0(\key_mem[5][46] ), .B1(n4273), .Y(
        n2459) );
  AO22X1 U1787 ( .A0(n4318), .A1(n674), .B0(\key_mem[3][46] ), .B1(n4338), .Y(
        n2203) );
  AO22X1 U1788 ( .A0(n3971), .A1(n1497), .B0(\key_mem[1][72] ), .B1(n3980), 
        .Y(n1921) );
  AO22X1 U1789 ( .A0(n3971), .A1(n1503), .B0(\key_mem[1][78] ), .B1(n3977), 
        .Y(n1915) );
  AO22X1 U1790 ( .A0(n4010), .A1(n1465), .B0(\key_mem[14][40] ), .B1(n4021), 
        .Y(n3617) );
  AO22X1 U1791 ( .A0(n4066), .A1(n1465), .B0(\key_mem[12][40] ), .B1(n4088), 
        .Y(n3361) );
  AO22X1 U1792 ( .A0(n4122), .A1(n1465), .B0(\key_mem[10][40] ), .B1(n4139), 
        .Y(n3105) );
  AO22X1 U1793 ( .A0(n4178), .A1(n1465), .B0(\key_mem[8][40] ), .B1(n4195), 
        .Y(n2849) );
  AO22X1 U1794 ( .A0(n4235), .A1(n1465), .B0(\key_mem[6][40] ), .B1(n4244), 
        .Y(n2593) );
  AO22X1 U1795 ( .A0(n4290), .A1(n1465), .B0(\key_mem[4][40] ), .B1(n4307), 
        .Y(n2337) );
  AO22X1 U1796 ( .A0(n4346), .A1(n1465), .B0(\key_mem[2][40] ), .B1(n4361), 
        .Y(n2081) );
  AO22X1 U1797 ( .A0(n3956), .A1(n1465), .B0(\key_mem[0][40] ), .B1(n1736), 
        .Y(n1825) );
  AO22X1 U1798 ( .A0(n4010), .A1(n1471), .B0(\key_mem[14][46] ), .B1(n4030), 
        .Y(n3611) );
  AO22X1 U1799 ( .A0(n4066), .A1(n1471), .B0(\key_mem[12][46] ), .B1(n4082), 
        .Y(n3355) );
  AO22X1 U1800 ( .A0(n4122), .A1(n1471), .B0(\key_mem[10][46] ), .B1(n4133), 
        .Y(n3099) );
  AO22X1 U1801 ( .A0(n4178), .A1(n1471), .B0(\key_mem[8][46] ), .B1(n4189), 
        .Y(n2843) );
  AO22X1 U1802 ( .A0(n4235), .A1(n1471), .B0(\key_mem[6][46] ), .B1(n4257), 
        .Y(n2587) );
  AO22X1 U1803 ( .A0(n4290), .A1(n1471), .B0(\key_mem[4][46] ), .B1(n4299), 
        .Y(n2331) );
  AO22X1 U1804 ( .A0(n4346), .A1(n1471), .B0(\key_mem[2][46] ), .B1(n4367), 
        .Y(n2075) );
  AO22X1 U1805 ( .A0(n3955), .A1(n1471), .B0(\key_mem[0][46] ), .B1(n3928), 
        .Y(n1819) );
  AO22X1 U1806 ( .A0(n4013), .A1(n1497), .B0(\key_mem[14][72] ), .B1(n4023), 
        .Y(n3585) );
  AO22X1 U1807 ( .A0(n4041), .A1(n1497), .B0(\key_mem[13][72] ), .B1(n4048), 
        .Y(n3457) );
  AO22X1 U1808 ( .A0(n4069), .A1(n1497), .B0(\key_mem[12][72] ), .B1(n4078), 
        .Y(n3329) );
  AO22X1 U1809 ( .A0(n4097), .A1(n1497), .B0(\key_mem[11][72] ), .B1(n4110), 
        .Y(n3201) );
  AO22X1 U1810 ( .A0(n4125), .A1(n1497), .B0(\key_mem[10][72] ), .B1(n4137), 
        .Y(n3073) );
  AO22X1 U1811 ( .A0(n4153), .A1(n1497), .B0(\key_mem[9][72] ), .B1(n4164), 
        .Y(n2945) );
  AO22X1 U1812 ( .A0(n4181), .A1(n648), .B0(\key_mem[8][72] ), .B1(n4195), .Y(
        n2817) );
  AO22X1 U1813 ( .A0(n4209), .A1(n1497), .B0(\key_mem[7][72] ), .B1(n4220), 
        .Y(n2689) );
  AO22X1 U1814 ( .A0(n4238), .A1(n648), .B0(\key_mem[6][72] ), .B1(n4244), .Y(
        n2561) );
  AO22X1 U1815 ( .A0(n4265), .A1(n1497), .B0(\key_mem[5][72] ), .B1(n4274), 
        .Y(n2433) );
  AO22X1 U1816 ( .A0(n4293), .A1(n648), .B0(\key_mem[4][72] ), .B1(n4306), .Y(
        n2305) );
  AO22X1 U1817 ( .A0(n4321), .A1(n1497), .B0(\key_mem[3][72] ), .B1(n4341), 
        .Y(n2177) );
  AO22X1 U1818 ( .A0(n4349), .A1(n648), .B0(\key_mem[2][72] ), .B1(n4369), .Y(
        n2049) );
  AO22X1 U1819 ( .A0(n3953), .A1(n648), .B0(\key_mem[0][72] ), .B1(n3931), .Y(
        n1793) );
  AO22X1 U1820 ( .A0(n4013), .A1(n1503), .B0(\key_mem[14][78] ), .B1(n4020), 
        .Y(n3579) );
  AO22X1 U1821 ( .A0(n4041), .A1(n1503), .B0(\key_mem[13][78] ), .B1(n4060), 
        .Y(n3451) );
  AO22X1 U1822 ( .A0(n4069), .A1(n1503), .B0(\key_mem[12][78] ), .B1(n4083), 
        .Y(n3323) );
  AO22X1 U1823 ( .A0(n4097), .A1(n1503), .B0(\key_mem[11][78] ), .B1(n4106), 
        .Y(n3195) );
  AO22X1 U1824 ( .A0(n4125), .A1(n1503), .B0(\key_mem[10][78] ), .B1(n4132), 
        .Y(n3067) );
  AO22X1 U1825 ( .A0(n4153), .A1(n1503), .B0(\key_mem[9][78] ), .B1(n4161), 
        .Y(n2939) );
  AO22X1 U1826 ( .A0(n4181), .A1(n642), .B0(\key_mem[8][78] ), .B1(n4188), .Y(
        n2811) );
  AO22X1 U1827 ( .A0(n4209), .A1(n1503), .B0(\key_mem[7][78] ), .B1(n4215), 
        .Y(n2683) );
  AO22X1 U1828 ( .A0(n4238), .A1(n642), .B0(\key_mem[6][78] ), .B1(n4248), .Y(
        n2555) );
  AO22X1 U1829 ( .A0(n4265), .A1(n1503), .B0(\key_mem[5][78] ), .B1(n4273), 
        .Y(n2427) );
  AO22X1 U1830 ( .A0(n4293), .A1(n642), .B0(\key_mem[4][78] ), .B1(n4306), .Y(
        n2299) );
  AO22X1 U1831 ( .A0(n4321), .A1(n1503), .B0(\key_mem[3][78] ), .B1(n4329), 
        .Y(n2171) );
  AO22X1 U1832 ( .A0(n4349), .A1(n642), .B0(\key_mem[2][78] ), .B1(n4366), .Y(
        n2043) );
  AO22X1 U1833 ( .A0(n3952), .A1(n642), .B0(\key_mem[0][78] ), .B1(n3931), .Y(
        n1787) );
  XNOR2X1 U1834 ( .A(n4882), .B(sboxw[8]), .Y(n9) );
  XNOR2X1 U1835 ( .A(n5079), .B(sboxw[14]), .Y(n10) );
  AOI222XL U1836 ( .A0(n1704), .A1(n795), .B0(key[115]), .B1(n1679), .C0(n1692), .C1(n796), .Y(n794) );
  INVX1 U1837 ( .A(n5224), .Y(n796) );
  OAI221XL U1838 ( .A0(n1665), .A1(n4824), .B0(n1659), .B1(n4823), .C0(n4822), 
        .Y(n3906) );
  INVX1 U1839 ( .A(key[6]), .Y(n4824) );
  INVX1 U1840 ( .A(n5736), .Y(n4823) );
  AOI221XL U1841 ( .A0(n1643), .A1(n53), .B0(n1624), .B1(key[134]), .C0(n4821), 
        .Y(n4822) );
  OAI221XL U1842 ( .A0(n1666), .A1(n4621), .B0(n1662), .B1(n4620), .C0(n4619), 
        .Y(n3880) );
  INVX1 U1843 ( .A(key[32]), .Y(n4621) );
  INVX1 U1844 ( .A(n5755), .Y(n4620) );
  AOI221XL U1845 ( .A0(n1648), .A1(n1127), .B0(n1622), .B1(key[160]), .C0(
        n4618), .Y(n4619) );
  OAI221XL U1846 ( .A0(n1665), .A1(n4812), .B0(n1662), .B1(n4811), .C0(n4810), 
        .Y(n3874) );
  INVX1 U1847 ( .A(key[38]), .Y(n4812) );
  INVX1 U1848 ( .A(n5737), .Y(n4811) );
  AOI221XL U1849 ( .A0(n1643), .A1(n1103), .B0(n1624), .B1(key[166]), .C0(
        n4809), .Y(n4810) );
  OAI221XL U1850 ( .A0(n1665), .A1(n4804), .B0(n1660), .B1(n4803), .C0(n4802), 
        .Y(n3842) );
  INVX1 U1851 ( .A(key[70]), .Y(n4804) );
  INVX1 U1852 ( .A(n5738), .Y(n4803) );
  AOI221XL U1853 ( .A0(n1643), .A1(n40), .B0(n1624), .B1(key[198]), .C0(n4801), 
        .Y(n4802) );
  OAI221XL U1854 ( .A0(n1666), .A1(n4608), .B0(n4607), .B1(n1655), .C0(n4606), 
        .Y(n3816) );
  INVX1 U1855 ( .A(key[96]), .Y(n4608) );
  AOI221XL U1856 ( .A0(n1636), .A1(n871), .B0(n1622), .B1(key[224]), .C0(n4605), .Y(n4606) );
  AO22X1 U1857 ( .A0(prev_key1_reg[96]), .A1(n1608), .B0(n1595), .B1(n4604), 
        .Y(n4605) );
  OAI221XL U1858 ( .A0(n1669), .A1(n5225), .B0(n5224), .B1(n1656), .C0(n5223), 
        .Y(n3797) );
  INVX1 U1859 ( .A(key[115]), .Y(n5225) );
  AOI221XL U1860 ( .A0(n1639), .A1(n795), .B0(n1627), .B1(key[243]), .C0(n5222), .Y(n5223) );
  AO22X1 U1861 ( .A0(prev_key1_reg[115]), .A1(n1611), .B0(n1598), .B1(n5221), 
        .Y(n5222) );
  OAI221XL U1862 ( .A0(n1676), .A1(n5086), .B0(n1652), .B1(n5085), .C0(n5084), 
        .Y(n3898) );
  INVX1 U1863 ( .A(key[14]), .Y(n5086) );
  INVX1 U1864 ( .A(n5713), .Y(n5085) );
  AOI221XL U1865 ( .A0(n1640), .A1(n10), .B0(n1625), .B1(key[142]), .C0(n5083), 
        .Y(n5084) );
  OAI221XL U1866 ( .A0(n1676), .A1(n5074), .B0(n1652), .B1(n5073), .C0(n5072), 
        .Y(n3866) );
  INVX1 U1867 ( .A(key[46]), .Y(n5074) );
  INVX1 U1868 ( .A(n5714), .Y(n5073) );
  AOI221XL U1869 ( .A0(n1641), .A1(n1071), .B0(n1625), .B1(key[174]), .C0(
        n5071), .Y(n5072) );
  XOR2X1 U1870 ( .A(n5088), .B(prev_key1_reg[111]), .Y(n5101) );
  XOR2X1 U1871 ( .A(n5286), .B(prev_key1_reg[117]), .Y(n5299) );
  XOR2X1 U1872 ( .A(n5351), .B(prev_key1_reg[119]), .Y(n5364) );
  XOR2X1 U1873 ( .A(n4858), .B(prev_key0_reg[104]), .Y(n4862) );
  XNOR2X1 U1874 ( .A(n4871), .B(prev_key1_reg[72]), .Y(n11) );
  OAI221XL U1875 ( .A0(n1667), .A1(n4889), .B0(n1660), .B1(n4888), .C0(n4887), 
        .Y(n3904) );
  INVX1 U1876 ( .A(key[8]), .Y(n4889) );
  INVX1 U1877 ( .A(n5730), .Y(n4888) );
  AOI221XL U1878 ( .A0(n1647), .A1(n9), .B0(n1634), .B1(key[136]), .C0(n4886), 
        .Y(n4887) );
  XOR3X1 U1879 ( .A(prev_key1_reg[47]), .B(prev_key1_reg[79]), .C(n5101), .Y(
        n5112) );
  XOR3X1 U1880 ( .A(prev_key1_reg[53]), .B(prev_key1_reg[85]), .C(n5299), .Y(
        n5310) );
  XOR3X1 U1881 ( .A(prev_key1_reg[55]), .B(prev_key1_reg[87]), .C(n5364), .Y(
        n5375) );
  AOI222XL U1882 ( .A0(n1716), .A1(n49), .B0(key[0]), .B1(n1685), .C0(n1700), 
        .C1(n5754), .Y(n1254) );
  AOI222XL U1883 ( .A0(n1705), .A1(n847), .B0(key[102]), .B1(n1680), .C0(n1693), .C1(n848), .Y(n846) );
  INVX1 U1884 ( .A(n1419), .Y(n845) );
  INVX1 U1885 ( .A(n4797), .Y(n848) );
  AOI222XL U1886 ( .A0(n1705), .A1(n839), .B0(key[104]), .B1(n1680), .C0(n1693), .C1(n840), .Y(n838) );
  INVX1 U1887 ( .A(n4862), .Y(n840) );
  AO22X1 U1888 ( .A0(n3964), .A1(n1425), .B0(\key_mem[1][0] ), .B1(n3984), .Y(
        n1993) );
  AO22X1 U1889 ( .A0(n3965), .A1(n1440), .B0(\key_mem[1][15] ), .B1(n3990), 
        .Y(n1978) );
  AO22X1 U1890 ( .A0(n3966), .A1(n1446), .B0(\key_mem[1][21] ), .B1(n3991), 
        .Y(n1972) );
  AO22X1 U1891 ( .A0(n3966), .A1(n1448), .B0(\key_mem[1][23] ), .B1(n3980), 
        .Y(n1970) );
  AO22X1 U1892 ( .A0(n3968), .A1(n1472), .B0(\key_mem[1][47] ), .B1(n3985), 
        .Y(n1946) );
  AO22X1 U1893 ( .A0(n3974), .A1(n1527), .B0(\key_mem[1][102] ), .B1(n3986), 
        .Y(n1891) );
  AO22X1 U1894 ( .A0(n3974), .A1(n1529), .B0(\key_mem[1][104] ), .B1(n3987), 
        .Y(n1889) );
  AO22X1 U1895 ( .A0(n4034), .A1(n1425), .B0(\key_mem[13][0] ), .B1(n4055), 
        .Y(n3529) );
  AO22X1 U1896 ( .A0(n4090), .A1(n720), .B0(\key_mem[11][0] ), .B1(n4117), .Y(
        n3273) );
  AO22X1 U1897 ( .A0(n4146), .A1(n720), .B0(\key_mem[9][0] ), .B1(n4173), .Y(
        n3017) );
  AO22X1 U1898 ( .A0(n4203), .A1(n720), .B0(\key_mem[7][0] ), .B1(n4214), .Y(
        n2761) );
  AO22X1 U1899 ( .A0(n4258), .A1(n720), .B0(\key_mem[5][0] ), .B1(n4283), .Y(
        n2505) );
  AO22X1 U1900 ( .A0(n4314), .A1(n720), .B0(\key_mem[3][0] ), .B1(n4337), .Y(
        n2249) );
  AO22X1 U1901 ( .A0(n4035), .A1(n1440), .B0(\key_mem[13][15] ), .B1(n4048), 
        .Y(n3514) );
  AO22X1 U1902 ( .A0(n4091), .A1(n705), .B0(\key_mem[11][15] ), .B1(n4104), 
        .Y(n3258) );
  AO22X1 U1903 ( .A0(n4147), .A1(n705), .B0(\key_mem[9][15] ), .B1(n735), .Y(
        n3002) );
  AO22X1 U1904 ( .A0(n4204), .A1(n705), .B0(\key_mem[7][15] ), .B1(n4221), .Y(
        n2746) );
  AO22X1 U1905 ( .A0(n4259), .A1(n705), .B0(\key_mem[5][15] ), .B1(n729), .Y(
        n2490) );
  AO22X1 U1906 ( .A0(n4315), .A1(n705), .B0(\key_mem[3][15] ), .B1(n4338), .Y(
        n2234) );
  AO22X1 U1907 ( .A0(n4036), .A1(n1446), .B0(\key_mem[13][21] ), .B1(n4049), 
        .Y(n3508) );
  AO22X1 U1908 ( .A0(n4092), .A1(n699), .B0(\key_mem[11][21] ), .B1(n4107), 
        .Y(n3252) );
  AO22X1 U1909 ( .A0(n4148), .A1(n699), .B0(\key_mem[9][21] ), .B1(n4171), .Y(
        n2996) );
  AO22X1 U1910 ( .A0(n4205), .A1(n699), .B0(\key_mem[7][21] ), .B1(n4221), .Y(
        n2740) );
  AO22X1 U1911 ( .A0(n4260), .A1(n699), .B0(\key_mem[5][21] ), .B1(n4283), .Y(
        n2484) );
  AO22X1 U1912 ( .A0(n4316), .A1(n699), .B0(\key_mem[3][21] ), .B1(n4338), .Y(
        n2228) );
  AO22X1 U1913 ( .A0(n4036), .A1(n1448), .B0(\key_mem[13][23] ), .B1(n4054), 
        .Y(n3506) );
  AO22X1 U1914 ( .A0(n4092), .A1(n697), .B0(\key_mem[11][23] ), .B1(n4107), 
        .Y(n3250) );
  AO22X1 U1915 ( .A0(n4148), .A1(n697), .B0(\key_mem[9][23] ), .B1(n4173), .Y(
        n2994) );
  AO22X1 U1916 ( .A0(n4205), .A1(n697), .B0(\key_mem[7][23] ), .B1(n4222), .Y(
        n2738) );
  AO22X1 U1917 ( .A0(n4260), .A1(n697), .B0(\key_mem[5][23] ), .B1(n4285), .Y(
        n2482) );
  AO22X1 U1918 ( .A0(n4316), .A1(n697), .B0(\key_mem[3][23] ), .B1(n4333), .Y(
        n2226) );
  AO22X1 U1919 ( .A0(n4038), .A1(n1472), .B0(\key_mem[13][47] ), .B1(n4061), 
        .Y(n3482) );
  AO22X1 U1920 ( .A0(n4094), .A1(n673), .B0(\key_mem[11][47] ), .B1(n4111), 
        .Y(n3226) );
  AO22X1 U1921 ( .A0(n4150), .A1(n673), .B0(\key_mem[9][47] ), .B1(n4171), .Y(
        n2970) );
  AO22X1 U1922 ( .A0(n732), .A1(n673), .B0(\key_mem[7][47] ), .B1(n4218), .Y(
        n2714) );
  AO22X1 U1923 ( .A0(n4262), .A1(n673), .B0(\key_mem[5][47] ), .B1(n4279), .Y(
        n2458) );
  AO22X1 U1924 ( .A0(n4318), .A1(n673), .B0(\key_mem[3][47] ), .B1(n4329), .Y(
        n2202) );
  AO22X1 U1925 ( .A0(n4044), .A1(n1527), .B0(\key_mem[13][102] ), .B1(n4057), 
        .Y(n3427) );
  AO22X1 U1926 ( .A0(n4100), .A1(n618), .B0(\key_mem[11][102] ), .B1(n4108), 
        .Y(n3171) );
  AO22X1 U1927 ( .A0(n4156), .A1(n618), .B0(\key_mem[9][102] ), .B1(n4170), 
        .Y(n2915) );
  AO22X1 U1928 ( .A0(n4212), .A1(n618), .B0(\key_mem[7][102] ), .B1(n4216), 
        .Y(n2659) );
  AO22X1 U1929 ( .A0(n4268), .A1(n618), .B0(\key_mem[5][102] ), .B1(n4282), 
        .Y(n2403) );
  AO22X1 U1930 ( .A0(n4324), .A1(n618), .B0(\key_mem[3][102] ), .B1(n4331), 
        .Y(n2147) );
  AO22X1 U1931 ( .A0(n4044), .A1(n1529), .B0(\key_mem[13][104] ), .B1(n4051), 
        .Y(n3425) );
  AO22X1 U1932 ( .A0(n4100), .A1(n616), .B0(\key_mem[11][104] ), .B1(n4105), 
        .Y(n3169) );
  AO22X1 U1933 ( .A0(n4156), .A1(n616), .B0(\key_mem[9][104] ), .B1(n4169), 
        .Y(n2913) );
  AO22X1 U1934 ( .A0(n4212), .A1(n616), .B0(\key_mem[7][104] ), .B1(n4224), 
        .Y(n2657) );
  AO22X1 U1935 ( .A0(n4268), .A1(n616), .B0(\key_mem[5][104] ), .B1(n4281), 
        .Y(n2401) );
  AO22X1 U1936 ( .A0(n4324), .A1(n616), .B0(\key_mem[3][104] ), .B1(n4336), 
        .Y(n2145) );
  AO22X1 U1937 ( .A0(n4006), .A1(n1425), .B0(\key_mem[14][0] ), .B1(n4023), 
        .Y(n3657) );
  AO22X1 U1938 ( .A0(n4062), .A1(n1425), .B0(\key_mem[12][0] ), .B1(n4088), 
        .Y(n3401) );
  AO22X1 U1939 ( .A0(n4118), .A1(n1425), .B0(\key_mem[10][0] ), .B1(n4139), 
        .Y(n3145) );
  AO22X1 U1940 ( .A0(n4174), .A1(n1425), .B0(\key_mem[8][0] ), .B1(n4195), .Y(
        n2889) );
  AO22X1 U1941 ( .A0(n4231), .A1(n1425), .B0(\key_mem[6][0] ), .B1(n4244), .Y(
        n2633) );
  AO22X1 U1942 ( .A0(n4286), .A1(n1425), .B0(\key_mem[4][0] ), .B1(n4302), .Y(
        n2377) );
  AO22X1 U1943 ( .A0(n4342), .A1(n1425), .B0(\key_mem[2][0] ), .B1(n4357), .Y(
        n2121) );
  AO22X1 U1944 ( .A0(n3960), .A1(n1425), .B0(\key_mem[0][0] ), .B1(n3930), .Y(
        n1865) );
  AO22X1 U1945 ( .A0(n4007), .A1(n1440), .B0(\key_mem[14][15] ), .B1(n4030), 
        .Y(n3642) );
  AO22X1 U1946 ( .A0(n4063), .A1(n1440), .B0(\key_mem[12][15] ), .B1(n4089), 
        .Y(n3386) );
  AO22X1 U1947 ( .A0(n4119), .A1(n1440), .B0(\key_mem[10][15] ), .B1(n736), 
        .Y(n3130) );
  AO22X1 U1948 ( .A0(n4175), .A1(n1440), .B0(\key_mem[8][15] ), .B1(n733), .Y(
        n2874) );
  AO22X1 U1949 ( .A0(n4232), .A1(n1440), .B0(\key_mem[6][15] ), .B1(n4249), 
        .Y(n2618) );
  AO22X1 U1950 ( .A0(n4287), .A1(n1440), .B0(\key_mem[4][15] ), .B1(n4305), 
        .Y(n2362) );
  AO22X1 U1951 ( .A0(n4343), .A1(n1440), .B0(\key_mem[2][15] ), .B1(n4360), 
        .Y(n2106) );
  AO22X1 U1952 ( .A0(n3958), .A1(n1440), .B0(\key_mem[0][15] ), .B1(n1720), 
        .Y(n1850) );
  AO22X1 U1953 ( .A0(n4008), .A1(n1446), .B0(\key_mem[14][21] ), .B1(n4031), 
        .Y(n3636) );
  AO22X1 U1954 ( .A0(n4064), .A1(n1446), .B0(\key_mem[12][21] ), .B1(n4086), 
        .Y(n3380) );
  AO22X1 U1955 ( .A0(n4120), .A1(n1446), .B0(\key_mem[10][21] ), .B1(n4143), 
        .Y(n3124) );
  AO22X1 U1956 ( .A0(n4176), .A1(n1446), .B0(\key_mem[8][21] ), .B1(n4199), 
        .Y(n2868) );
  AO22X1 U1957 ( .A0(n4233), .A1(n1446), .B0(\key_mem[6][21] ), .B1(n4248), 
        .Y(n2612) );
  AO22X1 U1958 ( .A0(n4288), .A1(n1446), .B0(\key_mem[4][21] ), .B1(n4305), 
        .Y(n2356) );
  AO22X1 U1959 ( .A0(n4344), .A1(n1446), .B0(\key_mem[2][21] ), .B1(n4357), 
        .Y(n2100) );
  AO22X1 U1960 ( .A0(n3958), .A1(n1446), .B0(\key_mem[0][21] ), .B1(n1728), 
        .Y(n1844) );
  AO22X1 U1961 ( .A0(n4008), .A1(n1448), .B0(\key_mem[14][23] ), .B1(n4024), 
        .Y(n3634) );
  AO22X1 U1962 ( .A0(n4064), .A1(n1448), .B0(\key_mem[12][23] ), .B1(n4089), 
        .Y(n3378) );
  AO22X1 U1963 ( .A0(n4120), .A1(n1448), .B0(\key_mem[10][23] ), .B1(n4145), 
        .Y(n3122) );
  AO22X1 U1964 ( .A0(n4176), .A1(n1448), .B0(\key_mem[8][23] ), .B1(n4201), 
        .Y(n2866) );
  AO22X1 U1965 ( .A0(n4233), .A1(n1448), .B0(\key_mem[6][23] ), .B1(n4256), 
        .Y(n2610) );
  AO22X1 U1966 ( .A0(n4288), .A1(n1448), .B0(\key_mem[4][23] ), .B1(n4310), 
        .Y(n2354) );
  AO22X1 U1967 ( .A0(n4344), .A1(n1448), .B0(\key_mem[2][23] ), .B1(n4355), 
        .Y(n2098) );
  AO22X1 U1968 ( .A0(n3957), .A1(n1448), .B0(\key_mem[0][23] ), .B1(n1728), 
        .Y(n1842) );
  AO22X1 U1969 ( .A0(n4010), .A1(n1472), .B0(\key_mem[14][47] ), .B1(n4032), 
        .Y(n3610) );
  AO22X1 U1970 ( .A0(n4066), .A1(n1472), .B0(\key_mem[12][47] ), .B1(n4081), 
        .Y(n3354) );
  AO22X1 U1971 ( .A0(n4122), .A1(n1472), .B0(\key_mem[10][47] ), .B1(n4145), 
        .Y(n3098) );
  AO22X1 U1972 ( .A0(n4178), .A1(n1472), .B0(\key_mem[8][47] ), .B1(n4201), 
        .Y(n2842) );
  AO22X1 U1973 ( .A0(n4235), .A1(n1472), .B0(\key_mem[6][47] ), .B1(n4257), 
        .Y(n2586) );
  AO22X1 U1974 ( .A0(n4290), .A1(n1472), .B0(\key_mem[4][47] ), .B1(n4311), 
        .Y(n2330) );
  AO22X1 U1975 ( .A0(n4346), .A1(n1472), .B0(\key_mem[2][47] ), .B1(n4368), 
        .Y(n2074) );
  AO22X1 U1976 ( .A0(n3955), .A1(n1472), .B0(\key_mem[0][47] ), .B1(n3928), 
        .Y(n1818) );
  AO22X1 U1977 ( .A0(n4016), .A1(n1527), .B0(\key_mem[14][102] ), .B1(n4026), 
        .Y(n3555) );
  AO22X1 U1978 ( .A0(n4072), .A1(n1527), .B0(\key_mem[12][102] ), .B1(n4087), 
        .Y(n3299) );
  AO22X1 U1979 ( .A0(n4128), .A1(n1527), .B0(\key_mem[10][102] ), .B1(n4141), 
        .Y(n3043) );
  AO22X1 U1980 ( .A0(n4184), .A1(n1527), .B0(\key_mem[8][102] ), .B1(n4197), 
        .Y(n2787) );
  AO22X1 U1981 ( .A0(n4241), .A1(n1527), .B0(\key_mem[6][102] ), .B1(n4253), 
        .Y(n2531) );
  AO22X1 U1982 ( .A0(n4296), .A1(n1527), .B0(\key_mem[4][102] ), .B1(n4306), 
        .Y(n2275) );
  AO22X1 U1983 ( .A0(n4352), .A1(n1527), .B0(\key_mem[2][102] ), .B1(n4364), 
        .Y(n2019) );
  AO22X1 U1984 ( .A0(n3950), .A1(n1527), .B0(\key_mem[0][102] ), .B1(n5761), 
        .Y(n1763) );
  AO22X1 U1985 ( .A0(n4016), .A1(n1529), .B0(\key_mem[14][104] ), .B1(n4027), 
        .Y(n3553) );
  AO22X1 U1986 ( .A0(n4072), .A1(n1529), .B0(\key_mem[12][104] ), .B1(n4084), 
        .Y(n3297) );
  AO22X1 U1987 ( .A0(n4128), .A1(n1529), .B0(\key_mem[10][104] ), .B1(n4141), 
        .Y(n3041) );
  AO22X1 U1988 ( .A0(n4184), .A1(n1529), .B0(\key_mem[8][104] ), .B1(n4197), 
        .Y(n2785) );
  AO22X1 U1989 ( .A0(n4241), .A1(n1529), .B0(\key_mem[6][104] ), .B1(n4248), 
        .Y(n2529) );
  AO22X1 U1990 ( .A0(n4296), .A1(n1529), .B0(\key_mem[4][104] ), .B1(n4309), 
        .Y(n2273) );
  AO22X1 U1991 ( .A0(n4352), .A1(n1529), .B0(\key_mem[2][104] ), .B1(n4356), 
        .Y(n2017) );
  AO22X1 U1992 ( .A0(n3949), .A1(n1529), .B0(\key_mem[0][104] ), .B1(n5761), 
        .Y(n1761) );
  XNOR2X1 U1993 ( .A(n5112), .B(sboxw[15]), .Y(n12) );
  XNOR2X1 U1994 ( .A(n5310), .B(sboxw[21]), .Y(n13) );
  XNOR2X1 U1995 ( .A(n5375), .B(sboxw[23]), .Y(n14) );
  AO22X1 U1996 ( .A0(sboxw[0]), .A1(n1608), .B0(n1595), .B1(n4629), .Y(n4630)
         );
  INVX1 U1997 ( .A(n1422), .Y(n4629) );
  OAI221XL U1998 ( .A0(n1667), .A1(n4877), .B0(n1661), .B1(n4876), .C0(n4875), 
        .Y(n3872) );
  INVX1 U1999 ( .A(key[40]), .Y(n4877) );
  AOI221XL U2000 ( .A0(n1647), .A1(n1095), .B0(n1633), .B1(key[168]), .C0(
        n4874), .Y(n4875) );
  INVX1 U2001 ( .A(n5731), .Y(n4876) );
  OAI221XL U2002 ( .A0(n1667), .A1(n4869), .B0(n1659), .B1(n4868), .C0(n4867), 
        .Y(n3840) );
  INVX1 U2003 ( .A(key[72]), .Y(n4869) );
  AOI221XL U2004 ( .A0(n1646), .A1(n11), .B0(n1633), .B1(key[200]), .C0(n4866), 
        .Y(n4867) );
  OAI221XL U2005 ( .A0(n1675), .A1(n5066), .B0(n1652), .B1(n4), .C0(n5065), 
        .Y(n3834) );
  AOI221XL U2006 ( .A0(n1641), .A1(n8), .B0(n1625), .B1(key[206]), .C0(n5064), 
        .Y(n5065) );
  OAI221XL U2007 ( .A0(n1675), .A1(n5061), .B0(n5060), .B1(n1657), .C0(n5059), 
        .Y(n3802) );
  INVX1 U2008 ( .A(key[110]), .Y(n5061) );
  AOI221XL U2009 ( .A0(n1641), .A1(n815), .B0(n1625), .B1(key[238]), .C0(n5058), .Y(n5059) );
  INVX1 U2010 ( .A(n5115), .Y(n1193) );
  AOI222XL U2011 ( .A0(n1713), .A1(n12), .B0(key[15]), .B1(n1689), .C0(n1699), 
        .C1(n5710), .Y(n1194) );
  INVX1 U2012 ( .A(n5313), .Y(n1169) );
  AOI222XL U2013 ( .A0(n1712), .A1(n13), .B0(key[21]), .B1(n1686), .C0(n1701), 
        .C1(n5692), .Y(n1170) );
  INVX1 U2014 ( .A(n5378), .Y(n1161) );
  AOI222XL U2015 ( .A0(n1712), .A1(n14), .B0(key[23]), .B1(n1685), .C0(n1703), 
        .C1(n5687), .Y(n1162) );
  INVX1 U2016 ( .A(n5103), .Y(n1065) );
  AOI222XL U2017 ( .A0(n1711), .A1(n1067), .B0(key[47]), .B1(n1684), .C0(n1698), .C1(n5711), .Y(n1066) );
  OAI221XL U2018 ( .A0(n1665), .A1(n4798), .B0(n4797), .B1(n1658), .C0(n4796), 
        .Y(n3810) );
  INVX1 U2019 ( .A(key[102]), .Y(n4798) );
  AOI221XL U2020 ( .A0(n1643), .A1(n847), .B0(n1624), .B1(key[230]), .C0(n4795), .Y(n4796) );
  AO22X1 U2021 ( .A0(prev_key1_reg[102]), .A1(n1619), .B0(n1606), .B1(n1419), 
        .Y(n4795) );
  OAI221XL U2022 ( .A0(n1667), .A1(n4863), .B0(n4862), .B1(n1658), .C0(n4861), 
        .Y(n3808) );
  INVX1 U2023 ( .A(key[104]), .Y(n4863) );
  AOI221XL U2024 ( .A0(n1648), .A1(n839), .B0(n1634), .B1(key[232]), .C0(n4860), .Y(n4861) );
  AO22X1 U2025 ( .A0(prev_key1_reg[104]), .A1(n1621), .B0(n1595), .B1(n4859), 
        .Y(n4860) );
  OAI221XL U2026 ( .A0(n1666), .A1(n4633), .B0(n1662), .B1(n4632), .C0(n4631), 
        .Y(n3912) );
  INVX1 U2027 ( .A(key[0]), .Y(n4633) );
  INVX1 U2028 ( .A(n5754), .Y(n4632) );
  AOI221XL U2029 ( .A0(n1644), .A1(n49), .B0(n1622), .B1(key[128]), .C0(n4630), 
        .Y(n4631) );
  XOR2X1 U2030 ( .A(n4891), .B(prev_key1_reg[105]), .Y(n4904) );
  INVX1 U2031 ( .A(n5169), .Y(n1057) );
  OAI221XL U2032 ( .A0(n1061), .A1(n4002), .B0(n3939), .B1(n5793), .C0(n1062), 
        .Y(n672) );
  INVX1 U2033 ( .A(n5136), .Y(n1061) );
  OAI221XL U2034 ( .A0(n1045), .A1(n3993), .B0(n3940), .B1(n5841), .C0(n1046), 
        .Y(n668) );
  INVX1 U2035 ( .A(n5268), .Y(n1045) );
  OAI221XL U2036 ( .A0(n933), .A1(n3996), .B0(n3943), .B1(n5795), .C0(n934), 
        .Y(n640) );
  INVX1 U2037 ( .A(n5128), .Y(n933) );
  OAI221XL U2038 ( .A0(n909), .A1(n3996), .B0(n3943), .B1(n5875), .C0(n910), 
        .Y(n634) );
  INVX1 U2039 ( .A(n5326), .Y(n909) );
  OAI221XL U2040 ( .A0(n1189), .A1(n4001), .B0(n3936), .B1(n5791), .C0(n1190), 
        .Y(n704) );
  INVX1 U2041 ( .A(n5148), .Y(n1189) );
  OAI221XL U2042 ( .A0(n1089), .A1(n4003), .B0(n3939), .B1(n5767), .C0(n1090), 
        .Y(n679) );
  INVX1 U2043 ( .A(n4906), .Y(n1089) );
  OAI221XL U2044 ( .A0(n1077), .A1(n4001), .B0(n3939), .B1(n5835), .C0(n1078), 
        .Y(n676) );
  OAI221XL U2045 ( .A0(n961), .A1(n3995), .B0(n3942), .B1(n5772), .C0(n962), 
        .Y(n647) );
  INVX1 U2046 ( .A(n4898), .Y(n961) );
  OAI221XL U2047 ( .A0(n949), .A1(n3995), .B0(n3942), .B1(n5833), .C0(n950), 
        .Y(n644) );
  XOR2X1 U2048 ( .A(n4990), .B(prev_key0_reg[108]), .Y(n4994) );
  XOR2X1 U2049 ( .A(n5121), .B(prev_key0_reg[112]), .Y(n5125) );
  XOR2X1 U2050 ( .A(n5253), .B(prev_key0_reg[116]), .Y(n5257) );
  XOR2X1 U2051 ( .A(new_sboxw[16]), .B(n295), .Y(n5411) );
  XOR2X1 U2052 ( .A(new_sboxw[19]), .B(n289), .Y(n5519) );
  XOR2X1 U2053 ( .A(new_sboxw[18]), .B(n291), .Y(n5483) );
  XOR2X1 U2054 ( .A(new_sboxw[20]), .B(n287), .Y(n5555) );
  XOR2X1 U2055 ( .A(new_sboxw[21]), .B(n285), .Y(n5591) );
  XOR2X1 U2056 ( .A(new_sboxw[22]), .B(n283), .Y(n5627) );
  XOR2X1 U2057 ( .A(n5383), .B(prev_key1_reg[96]), .Y(n4616) );
  XOR2X1 U2058 ( .A(n5455), .B(prev_key1_reg[98]), .Y(n4679) );
  XOR2X1 U2059 ( .A(n5491), .B(prev_key1_reg[99]), .Y(n4711) );
  XOR2X1 U2060 ( .A(n5563), .B(prev_key1_reg[101]), .Y(n4775) );
  XOR2X1 U2061 ( .A(n5599), .B(prev_key1_reg[102]), .Y(n4806) );
  XOR2X1 U2062 ( .A(n5635), .B(prev_key1_reg[103]), .Y(n4838) );
  XOR2X1 U2063 ( .A(n4924), .B(prev_key1_reg[106]), .Y(n4937) );
  XOR2X1 U2064 ( .A(n4957), .B(prev_key1_reg[107]), .Y(n4970) );
  XOR2X1 U2065 ( .A(n5023), .B(prev_key1_reg[109]), .Y(n5036) );
  XOR2X1 U2066 ( .A(n5527), .B(prev_key1_reg[100]), .Y(n4743) );
  XOR2X1 U2067 ( .A(n5121), .B(prev_key1_reg[112]), .Y(n5134) );
  XOR2X1 U2068 ( .A(n5154), .B(prev_key1_reg[113]), .Y(n5167) );
  XOR2X1 U2069 ( .A(n5187), .B(prev_key1_reg[114]), .Y(n5200) );
  XOR2X1 U2070 ( .A(n5253), .B(prev_key1_reg[116]), .Y(n5266) );
  XOR2X1 U2071 ( .A(n5319), .B(prev_key1_reg[118]), .Y(n5332) );
  XOR2X1 U2072 ( .A(n5419), .B(prev_key1_reg[97]), .Y(n4647) );
  XOR2X1 U2073 ( .A(n4990), .B(prev_key1_reg[108]), .Y(n5003) );
  INVX1 U2074 ( .A(n5161), .Y(n929) );
  OAI221XL U2075 ( .A0(n1205), .A1(n4002), .B0(n3936), .B1(n5837), .C0(n1206), 
        .Y(n708) );
  AOI222XL U2076 ( .A0(n1715), .A1(n33), .B0(key[12]), .B1(n1688), .C0(n1700), 
        .C1(n5718), .Y(n1206) );
  OAI221XL U2077 ( .A0(n1185), .A1(n4003), .B0(n3936), .B1(n5779), .C0(n1186), 
        .Y(n703) );
  INVX1 U2078 ( .A(n5181), .Y(n1185) );
  OAI221XL U2079 ( .A0(n1217), .A1(n4003), .B0(n3935), .B1(n5773), .C0(n1218), 
        .Y(n711) );
  INVX1 U2080 ( .A(n4918), .Y(n1217) );
  XOR2X1 U2081 ( .A(n5642), .B(prev_key0_reg[127]), .Y(n5685) );
  XOR2X1 U2082 ( .A(n5599), .B(prev_key0_reg[102]), .Y(n4797) );
  XOR2X1 U2083 ( .A(n5447), .B(prev_key0_reg[121]), .Y(n5423) );
  XOR2X1 U2084 ( .A(n5555), .B(prev_key0_reg[124]), .Y(n5531) );
  XOR2X1 U2085 ( .A(n5591), .B(prev_key0_reg[125]), .Y(n5567) );
  XOR2X1 U2086 ( .A(n5627), .B(prev_key0_reg[126]), .Y(n5603) );
  XOR2X1 U2087 ( .A(n5519), .B(prev_key0_reg[123]), .Y(n5495) );
  XOR2X1 U2088 ( .A(n5483), .B(prev_key0_reg[122]), .Y(n5459) );
  XOR2X1 U2089 ( .A(n5411), .B(prev_key0_reg[120]), .Y(n5387) );
  XOR2X1 U2090 ( .A(n5635), .B(prev_key0_reg[127]), .Y(n741) );
  XOR2X1 U2091 ( .A(n5383), .B(prev_key0_reg[96]), .Y(n4607) );
  XOR2X1 U2092 ( .A(n5419), .B(prev_key0_reg[97]), .Y(n4638) );
  XOR2X1 U2093 ( .A(n5491), .B(prev_key0_reg[99]), .Y(n4702) );
  XOR2X1 U2094 ( .A(n5527), .B(prev_key0_reg[100]), .Y(n4734) );
  XOR2X1 U2095 ( .A(n5563), .B(prev_key0_reg[101]), .Y(n4766) );
  XOR2X1 U2096 ( .A(n5635), .B(prev_key0_reg[103]), .Y(n4829) );
  XOR2X1 U2097 ( .A(n4924), .B(prev_key0_reg[106]), .Y(n4928) );
  XOR2X1 U2098 ( .A(n4957), .B(prev_key0_reg[107]), .Y(n4961) );
  XOR2X1 U2099 ( .A(n5023), .B(prev_key0_reg[109]), .Y(n5027) );
  XOR2X1 U2100 ( .A(n5088), .B(prev_key0_reg[111]), .Y(n5092) );
  XOR2X1 U2101 ( .A(n5154), .B(prev_key0_reg[113]), .Y(n5158) );
  XOR2X1 U2102 ( .A(n5187), .B(prev_key0_reg[114]), .Y(n5191) );
  XOR2X1 U2103 ( .A(n5286), .B(prev_key0_reg[117]), .Y(n5290) );
  XOR2X1 U2104 ( .A(n5319), .B(prev_key0_reg[118]), .Y(n5323) );
  XOR2X1 U2105 ( .A(n5351), .B(prev_key0_reg[119]), .Y(n5355) );
  XNOR2X1 U2106 ( .A(n4647), .B(prev_key1_reg[65]), .Y(n15) );
  XNOR2X1 U2107 ( .A(n4658), .B(sboxw[1]), .Y(n16) );
  INVX1 U2108 ( .A(n5260), .Y(n917) );
  AOI222XL U2109 ( .A0(n1707), .A1(n32), .B0(key[84]), .B1(n1682), .C0(n1695), 
        .C1(n5697), .Y(n918) );
  XOR3X1 U2110 ( .A(prev_key1_reg[35]), .B(prev_key1_reg[67]), .C(n4711), .Y(
        n4722) );
  XOR3X1 U2111 ( .A(prev_key1_reg[36]), .B(prev_key1_reg[68]), .C(n4743), .Y(
        n4754) );
  XOR3X1 U2112 ( .A(prev_key1_reg[37]), .B(prev_key1_reg[69]), .C(n4775), .Y(
        n4786) );
  XOR3X1 U2113 ( .A(prev_key1_reg[38]), .B(prev_key1_reg[70]), .C(n4806), .Y(
        n4817) );
  XOR3X1 U2114 ( .A(prev_key1_reg[39]), .B(prev_key1_reg[71]), .C(n4838), .Y(
        n4849) );
  XOR3X1 U2115 ( .A(prev_key1_reg[41]), .B(prev_key1_reg[73]), .C(n4904), .Y(
        n4915) );
  XOR3X1 U2116 ( .A(prev_key1_reg[42]), .B(prev_key1_reg[74]), .C(n4937), .Y(
        n4948) );
  XOR3X1 U2117 ( .A(prev_key1_reg[43]), .B(prev_key1_reg[75]), .C(n4970), .Y(
        n4981) );
  XOR3X1 U2118 ( .A(prev_key1_reg[45]), .B(prev_key1_reg[77]), .C(n5036), .Y(
        n5047) );
  XOR3X1 U2119 ( .A(prev_key1_reg[48]), .B(prev_key1_reg[80]), .C(n5134), .Y(
        n5145) );
  XOR3X1 U2120 ( .A(prev_key1_reg[49]), .B(prev_key1_reg[81]), .C(n5167), .Y(
        n5178) );
  XOR3X1 U2121 ( .A(prev_key1_reg[50]), .B(prev_key1_reg[82]), .C(n5200), .Y(
        n5211) );
  XOR3X1 U2122 ( .A(prev_key1_reg[52]), .B(prev_key1_reg[84]), .C(n5266), .Y(
        n5277) );
  XOR3X1 U2123 ( .A(prev_key1_reg[32]), .B(prev_key1_reg[64]), .C(n4616), .Y(
        n4626) );
  XOR3X1 U2124 ( .A(prev_key1_reg[33]), .B(prev_key1_reg[65]), .C(n4647), .Y(
        n4658) );
  XOR3X1 U2125 ( .A(prev_key1_reg[34]), .B(prev_key1_reg[66]), .C(n4679), .Y(
        n4690) );
  XOR3X1 U2126 ( .A(prev_key1_reg[44]), .B(prev_key1_reg[76]), .C(n5003), .Y(
        n5014) );
  XNOR3X1 U2127 ( .A(prev_key1_reg[57]), .B(n5435), .C(n5434), .Y(n17) );
  XNOR3X1 U2128 ( .A(prev_key1_reg[60]), .B(n5543), .C(n5542), .Y(n18) );
  XNOR3X1 U2129 ( .A(prev_key1_reg[61]), .B(n5579), .C(n5578), .Y(n19) );
  XNOR3X1 U2130 ( .A(prev_key1_reg[62]), .B(n5615), .C(n5614), .Y(n20) );
  XNOR3X1 U2131 ( .A(prev_key1_reg[59]), .B(n5507), .C(n5506), .Y(n21) );
  XNOR3X1 U2132 ( .A(prev_key1_reg[58]), .B(n5471), .C(n5470), .Y(n22) );
  XNOR3X1 U2133 ( .A(prev_key1_reg[56]), .B(n5399), .C(n5398), .Y(n23) );
  XNOR3X1 U2134 ( .A(sboxw[25]), .B(prev_key1_reg[57]), .C(n5448), .Y(n24) );
  XNOR3X1 U2135 ( .A(sboxw[28]), .B(prev_key1_reg[60]), .C(n5556), .Y(n25) );
  XNOR3X1 U2136 ( .A(sboxw[29]), .B(prev_key1_reg[61]), .C(n5592), .Y(n26) );
  XNOR3X1 U2137 ( .A(sboxw[30]), .B(prev_key1_reg[62]), .C(n5628), .Y(n27) );
  XNOR3X1 U2138 ( .A(sboxw[27]), .B(prev_key1_reg[59]), .C(n5520), .Y(n28) );
  XNOR3X1 U2139 ( .A(sboxw[26]), .B(prev_key1_reg[58]), .C(n5484), .Y(n29) );
  XNOR3X1 U2140 ( .A(sboxw[24]), .B(prev_key1_reg[56]), .C(n5412), .Y(n30) );
  XOR2X1 U2141 ( .A(n5642), .B(prev_key1_reg[127]), .Y(n5686) );
  XOR3X1 U2142 ( .A(prev_key1_reg[54]), .B(prev_key1_reg[86]), .C(n5332), .Y(
        n5342) );
  AOI222XL U2143 ( .A0(n1712), .A1(n24), .B0(key[25]), .B1(n1690), .C0(n1700), 
        .C1(n1156), .Y(n1154) );
  INVX1 U2144 ( .A(n5453), .Y(n1156) );
  AOI222XL U2145 ( .A0(n1710), .A1(n17), .B0(key[57]), .B1(n1683), .C0(n1697), 
        .C1(n1028), .Y(n1026) );
  INVX1 U2146 ( .A(n5440), .Y(n1028) );
  AOI222XL U2147 ( .A0(n1706), .A1(n899), .B0(key[89]), .B1(n1681), .C0(n1694), 
        .C1(n900), .Y(n898) );
  INVX1 U2148 ( .A(n5430), .Y(n900) );
  AOI222XL U2149 ( .A0(n1716), .A1(n59), .B0(key[121]), .B1(n1678), .C0(n1691), 
        .C1(n772), .Y(n770) );
  INVX1 U2150 ( .A(n5423), .Y(n772) );
  AOI222XL U2151 ( .A0(n1712), .A1(n25), .B0(key[28]), .B1(n1686), .C0(n1703), 
        .C1(n1144), .Y(n1142) );
  INVX1 U2152 ( .A(n5561), .Y(n1144) );
  AOI222XL U2153 ( .A0(n1709), .A1(n18), .B0(key[60]), .B1(n1687), .C0(n1696), 
        .C1(n1016), .Y(n1014) );
  INVX1 U2154 ( .A(n5548), .Y(n1016) );
  AOI222XL U2155 ( .A0(n1706), .A1(n887), .B0(key[92]), .B1(n1681), .C0(n1694), 
        .C1(n888), .Y(n886) );
  INVX1 U2156 ( .A(n5538), .Y(n888) );
  AOI222XL U2157 ( .A0(n1715), .A1(n60), .B0(key[124]), .B1(n1678), .C0(n1691), 
        .C1(n760), .Y(n758) );
  INVX1 U2158 ( .A(n5531), .Y(n760) );
  AOI222XL U2159 ( .A0(n1716), .A1(n26), .B0(key[29]), .B1(n1686), .C0(n1701), 
        .C1(n1140), .Y(n1138) );
  INVX1 U2160 ( .A(n5597), .Y(n1140) );
  AOI222XL U2161 ( .A0(n1709), .A1(n19), .B0(key[61]), .B1(n1688), .C0(n1696), 
        .C1(n1012), .Y(n1010) );
  INVX1 U2162 ( .A(n5584), .Y(n1012) );
  AOI222XL U2163 ( .A0(n1706), .A1(n883), .B0(key[93]), .B1(n1681), .C0(n1694), 
        .C1(n884), .Y(n882) );
  INVX1 U2164 ( .A(n5574), .Y(n884) );
  AOI222XL U2165 ( .A0(n5759), .A1(n61), .B0(key[125]), .B1(n1678), .C0(n1691), 
        .C1(n756), .Y(n754) );
  INVX1 U2166 ( .A(n5567), .Y(n756) );
  AOI222XL U2167 ( .A0(n1713), .A1(n27), .B0(key[30]), .B1(n1686), .C0(n1700), 
        .C1(n1136), .Y(n1134) );
  INVX1 U2168 ( .A(n5633), .Y(n1136) );
  AOI222XL U2169 ( .A0(n1709), .A1(n20), .B0(key[62]), .B1(n1689), .C0(n1696), 
        .C1(n1008), .Y(n1006) );
  INVX1 U2170 ( .A(n5620), .Y(n1008) );
  AOI222XL U2171 ( .A0(n1706), .A1(n879), .B0(key[94]), .B1(n1681), .C0(n1694), 
        .C1(n880), .Y(n878) );
  INVX1 U2172 ( .A(n5610), .Y(n880) );
  AOI222XL U2173 ( .A0(n1714), .A1(n62), .B0(key[126]), .B1(n1678), .C0(n1691), 
        .C1(n752), .Y(n750) );
  INVX1 U2174 ( .A(n5603), .Y(n752) );
  AOI222XL U2175 ( .A0(n1712), .A1(n28), .B0(key[27]), .B1(n5757), .C0(n1699), 
        .C1(n1148), .Y(n1146) );
  INVX1 U2176 ( .A(n5525), .Y(n1148) );
  AOI222XL U2177 ( .A0(n1709), .A1(n21), .B0(key[59]), .B1(n1688), .C0(n1696), 
        .C1(n1020), .Y(n1018) );
  INVX1 U2178 ( .A(n5512), .Y(n1020) );
  AOI222XL U2179 ( .A0(n1706), .A1(n891), .B0(key[91]), .B1(n1681), .C0(n1694), 
        .C1(n892), .Y(n890) );
  INVX1 U2180 ( .A(n5502), .Y(n892) );
  AOI222XL U2181 ( .A0(n1715), .A1(n63), .B0(key[123]), .B1(n1678), .C0(n1691), 
        .C1(n764), .Y(n762) );
  INVX1 U2182 ( .A(n5495), .Y(n764) );
  AOI222XL U2183 ( .A0(n1712), .A1(n29), .B0(key[26]), .B1(n1688), .C0(n5758), 
        .C1(n1152), .Y(n1150) );
  INVX1 U2184 ( .A(n5489), .Y(n1152) );
  AOI222XL U2185 ( .A0(n1710), .A1(n22), .B0(key[58]), .B1(n1690), .C0(n1697), 
        .C1(n1024), .Y(n1022) );
  INVX1 U2186 ( .A(n5476), .Y(n1024) );
  AOI222XL U2187 ( .A0(n1706), .A1(n895), .B0(key[90]), .B1(n1681), .C0(n1694), 
        .C1(n896), .Y(n894) );
  INVX1 U2188 ( .A(n5466), .Y(n896) );
  AOI222XL U2189 ( .A0(n1716), .A1(n64), .B0(key[122]), .B1(n1678), .C0(n1691), 
        .C1(n768), .Y(n766) );
  INVX1 U2190 ( .A(n5459), .Y(n768) );
  AOI222XL U2191 ( .A0(n1712), .A1(n30), .B0(key[24]), .B1(n5757), .C0(n1701), 
        .C1(n1160), .Y(n1158) );
  INVX1 U2192 ( .A(n5417), .Y(n1160) );
  AOI222XL U2193 ( .A0(n1710), .A1(n23), .B0(key[56]), .B1(n1683), .C0(n1697), 
        .C1(n1032), .Y(n1030) );
  INVX1 U2194 ( .A(n5404), .Y(n1032) );
  AOI222XL U2195 ( .A0(n1707), .A1(n903), .B0(key[88]), .B1(n1681), .C0(n1700), 
        .C1(n904), .Y(n902) );
  INVX1 U2196 ( .A(n5394), .Y(n904) );
  AOI222XL U2197 ( .A0(n1713), .A1(n65), .B0(key[120]), .B1(n1678), .C0(n1691), 
        .C1(n776), .Y(n774) );
  INVX1 U2198 ( .A(n5387), .Y(n776) );
  AOI222XL U2199 ( .A0(n1706), .A1(n5684), .B0(key[95]), .B1(n1681), .C0(n1694), .C1(n5683), .Y(n874) );
  AOI222XL U2200 ( .A0(n5759), .A1(n5686), .B0(key[127]), .B1(n1678), .C0(
        n1691), .C1(n5685), .Y(n743) );
  INVX1 U2201 ( .A(n4693), .Y(n1245) );
  AOI222XL U2202 ( .A0(n1715), .A1(n50), .B0(key[2]), .B1(n1685), .C0(n1702), 
        .C1(n5748), .Y(n1246) );
  INVX1 U2203 ( .A(n4725), .Y(n1241) );
  AOI222XL U2204 ( .A0(n1714), .A1(n51), .B0(key[3]), .B1(n1689), .C0(n1703), 
        .C1(n5745), .Y(n1242) );
  INVX1 U2205 ( .A(n4789), .Y(n1233) );
  AOI222XL U2206 ( .A0(n1716), .A1(n52), .B0(key[5]), .B1(n1690), .C0(n1701), 
        .C1(n5739), .Y(n1234) );
  INVX1 U2207 ( .A(n4852), .Y(n1225) );
  AOI222XL U2208 ( .A0(n1715), .A1(n54), .B0(key[7]), .B1(n1687), .C0(n1699), 
        .C1(n5733), .Y(n1226) );
  INVX1 U2209 ( .A(n5345), .Y(n1165) );
  INVX1 U2210 ( .A(n4681), .Y(n1117) );
  AOI222XL U2211 ( .A0(n1713), .A1(n1119), .B0(key[34]), .B1(n1686), .C0(n1700), .C1(n5749), .Y(n1118) );
  INVX1 U2212 ( .A(n4713), .Y(n1113) );
  AOI222XL U2213 ( .A0(n5759), .A1(n1115), .B0(key[35]), .B1(n1685), .C0(n1702), .C1(n5746), .Y(n1114) );
  INVX1 U2214 ( .A(n4777), .Y(n1105) );
  AOI222XL U2215 ( .A0(n1710), .A1(n1107), .B0(key[37]), .B1(n1686), .C0(n1703), .C1(n5740), .Y(n1106) );
  INVX1 U2216 ( .A(n4840), .Y(n1097) );
  AOI222XL U2217 ( .A0(n1711), .A1(n1099), .B0(key[39]), .B1(n1684), .C0(n1698), .C1(n5734), .Y(n1098) );
  AOI222XL U2218 ( .A0(n1709), .A1(n37), .B0(key[66]), .B1(n1690), .C0(n1696), 
        .C1(n5750), .Y(n990) );
  INVX1 U2219 ( .A(n4673), .Y(n989) );
  AOI222XL U2220 ( .A0(n1709), .A1(n38), .B0(key[67]), .B1(n1687), .C0(n1696), 
        .C1(n5747), .Y(n986) );
  INVX1 U2221 ( .A(n4705), .Y(n985) );
  AOI222XL U2222 ( .A0(n1708), .A1(n39), .B0(key[69]), .B1(n1689), .C0(n1695), 
        .C1(n5741), .Y(n978) );
  INVX1 U2223 ( .A(n4769), .Y(n977) );
  AOI222XL U2224 ( .A0(n1708), .A1(n41), .B0(key[71]), .B1(n1688), .C0(n1695), 
        .C1(n5735), .Y(n970) );
  INVX1 U2225 ( .A(n4832), .Y(n969) );
  AOI222XL U2226 ( .A0(n1706), .A1(n867), .B0(key[97]), .B1(n1681), .C0(n1694), 
        .C1(n868), .Y(n866) );
  INVX1 U2227 ( .A(n4638), .Y(n868) );
  AOI222XL U2228 ( .A0(n1706), .A1(n863), .B0(key[98]), .B1(n1680), .C0(n1694), 
        .C1(n864), .Y(n862) );
  INVX1 U2229 ( .A(n4670), .Y(n864) );
  AOI222XL U2230 ( .A0(n1705), .A1(n859), .B0(key[99]), .B1(n1680), .C0(n1693), 
        .C1(n860), .Y(n858) );
  INVX1 U2231 ( .A(n4702), .Y(n860) );
  AOI222XL U2232 ( .A0(n1705), .A1(n855), .B0(key[100]), .B1(n1680), .C0(n1693), .C1(n856), .Y(n854) );
  INVX1 U2233 ( .A(n4734), .Y(n856) );
  AOI222XL U2234 ( .A0(n1705), .A1(n851), .B0(key[101]), .B1(n1680), .C0(n1693), .C1(n852), .Y(n850) );
  INVX1 U2235 ( .A(n4766), .Y(n852) );
  AOI222XL U2236 ( .A0(n1705), .A1(n843), .B0(key[103]), .B1(n1680), .C0(n1693), .C1(n844), .Y(n842) );
  INVX1 U2237 ( .A(n4829), .Y(n844) );
  AOI222XL U2238 ( .A0(n1705), .A1(n831), .B0(key[106]), .B1(n1680), .C0(n1693), .C1(n832), .Y(n830) );
  INVX1 U2239 ( .A(n4928), .Y(n832) );
  AOI222XL U2240 ( .A0(n1705), .A1(n823), .B0(key[108]), .B1(n1679), .C0(n1693), .C1(n824), .Y(n822) );
  INVX1 U2241 ( .A(n4994), .Y(n824) );
  AOI222XL U2242 ( .A0(n1704), .A1(n819), .B0(key[109]), .B1(n1679), .C0(n1692), .C1(n820), .Y(n818) );
  INVX1 U2243 ( .A(n5027), .Y(n820) );
  AOI222XL U2244 ( .A0(n1704), .A1(n811), .B0(key[111]), .B1(n1679), .C0(n1692), .C1(n812), .Y(n810) );
  INVX1 U2245 ( .A(n5092), .Y(n812) );
  AOI222XL U2246 ( .A0(n1704), .A1(n807), .B0(key[112]), .B1(n1679), .C0(n1692), .C1(n808), .Y(n806) );
  INVX1 U2247 ( .A(n5125), .Y(n808) );
  AOI222XL U2248 ( .A0(n1704), .A1(n803), .B0(key[113]), .B1(n1679), .C0(n1692), .C1(n804), .Y(n802) );
  INVX1 U2249 ( .A(n5158), .Y(n804) );
  AOI222XL U2250 ( .A0(n1704), .A1(n799), .B0(key[114]), .B1(n1679), .C0(n1692), .C1(n800), .Y(n798) );
  INVX1 U2251 ( .A(n5191), .Y(n800) );
  AOI222XL U2252 ( .A0(n1704), .A1(n791), .B0(key[116]), .B1(n1679), .C0(n1692), .C1(n792), .Y(n790) );
  INVX1 U2253 ( .A(n5257), .Y(n792) );
  AOI222XL U2254 ( .A0(n1704), .A1(n787), .B0(key[117]), .B1(n1679), .C0(n1692), .C1(n788), .Y(n786) );
  INVX1 U2255 ( .A(n5290), .Y(n788) );
  AOI222XL U2256 ( .A0(n1704), .A1(n783), .B0(key[118]), .B1(n1678), .C0(n1692), .C1(n784), .Y(n782) );
  INVX1 U2257 ( .A(n5323), .Y(n784) );
  AOI222XL U2258 ( .A0(n5759), .A1(n779), .B0(key[119]), .B1(n1678), .C0(n1691), .C1(n780), .Y(n778) );
  INVX1 U2259 ( .A(n5355), .Y(n780) );
  XOR3X1 U2260 ( .A(prev_key1_reg[63]), .B(n5665), .C(n5651), .Y(n5682) );
  XOR3X1 U2261 ( .A(sboxw[31]), .B(prev_key1_reg[63]), .C(n5684), .Y(n5680) );
  OAI221XL U2262 ( .A0(n1173), .A1(n4004), .B0(n3937), .B1(n5839), .C0(n1174), 
        .Y(n700) );
  INVX1 U2263 ( .A(n5280), .Y(n1173) );
  AO22X1 U2264 ( .A0(sboxw[1]), .A1(n1608), .B0(n1595), .B1(n4661), .Y(n4662)
         );
  AO22X1 U2265 ( .A0(prev_key1_reg[33]), .A1(n1608), .B0(n1595), .B1(n4649), 
        .Y(n4650) );
  AO22X1 U2266 ( .A0(prev_key1_reg[65]), .A1(n1608), .B0(n1595), .B1(n4641), 
        .Y(n4642) );
  XOR2X1 U2267 ( .A(new_sboxw[23]), .B(rcon_reg[7]), .Y(n5642) );
  AO22X1 U2268 ( .A0(sboxw[2]), .A1(n1618), .B0(n1606), .B1(n4693), .Y(n4694)
         );
  AO22X1 U2269 ( .A0(sboxw[3]), .A1(n1621), .B0(n1603), .B1(n4725), .Y(n4726)
         );
  AO22X1 U2270 ( .A0(sboxw[5]), .A1(n1619), .B0(n1606), .B1(n4789), .Y(n4790)
         );
  AO22X1 U2271 ( .A0(sboxw[7]), .A1(n1616), .B0(n1607), .B1(n4852), .Y(n4853)
         );
  AO22X1 U2272 ( .A0(sboxw[10]), .A1(n1621), .B0(n1605), .B1(n4951), .Y(n4952)
         );
  AO22X1 U2273 ( .A0(sboxw[13]), .A1(n1609), .B0(n1596), .B1(n5050), .Y(n5051)
         );
  AO22X1 U2274 ( .A0(sboxw[15]), .A1(n1610), .B0(n1597), .B1(n5115), .Y(n5116)
         );
  AO22X1 U2275 ( .A0(prev_key1_reg[34]), .A1(n1619), .B0(n1602), .B1(n4681), 
        .Y(n4682) );
  AO22X1 U2276 ( .A0(prev_key1_reg[35]), .A1(n1620), .B0(n1605), .B1(n4713), 
        .Y(n4714) );
  AO22X1 U2277 ( .A0(prev_key1_reg[37]), .A1(n1617), .B0(n1603), .B1(n4777), 
        .Y(n4778) );
  AO22X1 U2278 ( .A0(prev_key1_reg[39]), .A1(n1620), .B0(n1607), .B1(n4840), 
        .Y(n4841) );
  AO22X1 U2279 ( .A0(prev_key1_reg[42]), .A1(n1618), .B0(n1606), .B1(n4939), 
        .Y(n4940) );
  AO22X1 U2280 ( .A0(prev_key1_reg[45]), .A1(n1609), .B0(n1596), .B1(n5038), 
        .Y(n5039) );
  AO22X1 U2281 ( .A0(prev_key1_reg[47]), .A1(n1610), .B0(n1597), .B1(n5103), 
        .Y(n5104) );
  AO22X1 U2282 ( .A0(prev_key1_reg[66]), .A1(n1608), .B0(n1595), .B1(n4673), 
        .Y(n4674) );
  AO22X1 U2283 ( .A0(prev_key1_reg[67]), .A1(n1621), .B0(n1604), .B1(n4705), 
        .Y(n4706) );
  AO22X1 U2284 ( .A0(prev_key1_reg[69]), .A1(n1620), .B0(n1602), .B1(n4769), 
        .Y(n4770) );
  AO22X1 U2285 ( .A0(prev_key1_reg[71]), .A1(n1621), .B0(n1605), .B1(n4832), 
        .Y(n4833) );
  AO22X1 U2286 ( .A0(prev_key1_reg[74]), .A1(n1617), .B0(n1604), .B1(n4931), 
        .Y(n4932) );
  AO22X1 U2287 ( .A0(prev_key1_reg[77]), .A1(n1609), .B0(n1596), .B1(n5030), 
        .Y(n5031) );
  AO22X1 U2288 ( .A0(prev_key1_reg[79]), .A1(n1610), .B0(n1597), .B1(n5095), 
        .Y(n5096) );
  AO22X1 U2289 ( .A0(sboxw[9]), .A1(n1621), .B0(n5668), .B1(n4918), .Y(n4919)
         );
  AO22X1 U2290 ( .A0(prev_key1_reg[41]), .A1(n1621), .B0(n5668), .B1(n4906), 
        .Y(n4907) );
  AO22X1 U2291 ( .A0(prev_key1_reg[73]), .A1(n1616), .B0(n1603), .B1(n4898), 
        .Y(n4899) );
  AO22X1 U2292 ( .A0(sboxw[14]), .A1(n1609), .B0(n1596), .B1(n5082), .Y(n5083)
         );
  AO22X1 U2293 ( .A0(prev_key1_reg[46]), .A1(n1609), .B0(n1596), .B1(n5070), 
        .Y(n5071) );
  AO22X1 U2294 ( .A0(prev_key1_reg[36]), .A1(n1621), .B0(n1603), .B1(n4745), 
        .Y(n4746) );
  XNOR2X1 U2295 ( .A(n4904), .B(prev_key1_reg[73]), .Y(n31) );
  AO22X1 U2296 ( .A0(sboxw[20]), .A1(n1612), .B0(n1599), .B1(n5280), .Y(n5281)
         );
  AO22X1 U2297 ( .A0(prev_key1_reg[52]), .A1(n1612), .B0(n1599), .B1(n5268), 
        .Y(n5269) );
  AO22X1 U2298 ( .A0(prev_key1_reg[84]), .A1(n1612), .B0(n1599), .B1(n5260), 
        .Y(n5261) );
  AO22X1 U2299 ( .A0(n3964), .A1(n1426), .B0(\key_mem[1][1] ), .B1(n3984), .Y(
        n1992) );
  AO22X1 U2300 ( .A0(n3964), .A1(n1427), .B0(\key_mem[1][2] ), .B1(n3982), .Y(
        n1991) );
  AO22X1 U2301 ( .A0(n3964), .A1(n1428), .B0(\key_mem[1][3] ), .B1(n3981), .Y(
        n1990) );
  AO22X1 U2302 ( .A0(n3964), .A1(n1429), .B0(\key_mem[1][4] ), .B1(n3980), .Y(
        n1989) );
  AO22X1 U2303 ( .A0(n3964), .A1(n1430), .B0(\key_mem[1][5] ), .B1(n3984), .Y(
        n1988) );
  AO22X1 U2304 ( .A0(n3964), .A1(n1432), .B0(\key_mem[1][7] ), .B1(n3985), .Y(
        n1986) );
  AO22X1 U2305 ( .A0(n3965), .A1(n1435), .B0(\key_mem[1][10] ), .B1(n3990), 
        .Y(n1983) );
  AO22X1 U2306 ( .A0(n3965), .A1(n1438), .B0(\key_mem[1][13] ), .B1(n3991), 
        .Y(n1980) );
  AO22X1 U2307 ( .A0(n3965), .A1(n1443), .B0(\key_mem[1][18] ), .B1(n3988), 
        .Y(n1975) );
  AO22X1 U2308 ( .A0(n3966), .A1(n1447), .B0(\key_mem[1][22] ), .B1(n3987), 
        .Y(n1971) );
  AO22X1 U2309 ( .A0(n3966), .A1(n1449), .B0(\key_mem[1][24] ), .B1(n3990), 
        .Y(n1969) );
  AO22X1 U2310 ( .A0(n3966), .A1(n1450), .B0(\key_mem[1][25] ), .B1(n3988), 
        .Y(n1968) );
  AO22X1 U2311 ( .A0(n3966), .A1(n1451), .B0(\key_mem[1][26] ), .B1(n3978), 
        .Y(n1967) );
  AO22X1 U2312 ( .A0(n3966), .A1(n1452), .B0(\key_mem[1][27] ), .B1(n3989), 
        .Y(n1966) );
  AO22X1 U2313 ( .A0(n3966), .A1(n1453), .B0(\key_mem[1][28] ), .B1(n3990), 
        .Y(n1965) );
  AO22X1 U2314 ( .A0(n3966), .A1(n1454), .B0(\key_mem[1][29] ), .B1(n3991), 
        .Y(n1964) );
  AO22X1 U2315 ( .A0(n3967), .A1(n1455), .B0(\key_mem[1][30] ), .B1(n3991), 
        .Y(n1963) );
  AO22X1 U2316 ( .A0(n3967), .A1(n1456), .B0(\key_mem[1][31] ), .B1(n3986), 
        .Y(n1962) );
  AO22X1 U2317 ( .A0(n3967), .A1(n1458), .B0(\key_mem[1][33] ), .B1(n3977), 
        .Y(n1960) );
  AO22X1 U2318 ( .A0(n3967), .A1(n1459), .B0(\key_mem[1][34] ), .B1(n3989), 
        .Y(n1959) );
  AO22X1 U2319 ( .A0(n3967), .A1(n1460), .B0(\key_mem[1][35] ), .B1(n3986), 
        .Y(n1958) );
  AO22X1 U2320 ( .A0(n3967), .A1(n1461), .B0(\key_mem[1][36] ), .B1(n3988), 
        .Y(n1957) );
  AO22X1 U2321 ( .A0(n3967), .A1(n1462), .B0(\key_mem[1][37] ), .B1(n3989), 
        .Y(n1956) );
  AO22X1 U2322 ( .A0(n3967), .A1(n1464), .B0(\key_mem[1][39] ), .B1(n3987), 
        .Y(n1954) );
  AO22X1 U2323 ( .A0(n3968), .A1(n1467), .B0(\key_mem[1][42] ), .B1(n3986), 
        .Y(n1951) );
  AO22X1 U2324 ( .A0(n3968), .A1(n1470), .B0(\key_mem[1][45] ), .B1(n3989), 
        .Y(n1948) );
  AO22X1 U2325 ( .A0(n3969), .A1(n1475), .B0(\key_mem[1][50] ), .B1(n3989), 
        .Y(n1943) );
  AO22X1 U2326 ( .A0(n3969), .A1(n1478), .B0(\key_mem[1][53] ), .B1(n3989), 
        .Y(n1940) );
  AO22X1 U2327 ( .A0(n3969), .A1(n1480), .B0(\key_mem[1][55] ), .B1(n3986), 
        .Y(n1938) );
  AO22X1 U2328 ( .A0(n3969), .A1(n1481), .B0(\key_mem[1][56] ), .B1(n3981), 
        .Y(n1937) );
  AO22X1 U2329 ( .A0(n3969), .A1(n1482), .B0(\key_mem[1][57] ), .B1(n3980), 
        .Y(n1936) );
  AO22X1 U2330 ( .A0(n3969), .A1(n1483), .B0(\key_mem[1][58] ), .B1(n3979), 
        .Y(n1935) );
  AO22X1 U2331 ( .A0(n3969), .A1(n1484), .B0(\key_mem[1][59] ), .B1(n3978), 
        .Y(n1934) );
  AO22X1 U2332 ( .A0(n3970), .A1(n1485), .B0(\key_mem[1][60] ), .B1(n3977), 
        .Y(n1933) );
  AO22X1 U2333 ( .A0(n3970), .A1(n1486), .B0(\key_mem[1][61] ), .B1(n3981), 
        .Y(n1932) );
  AO22X1 U2334 ( .A0(n3970), .A1(n1487), .B0(\key_mem[1][62] ), .B1(n3980), 
        .Y(n1931) );
  AO22X1 U2335 ( .A0(n3970), .A1(n1488), .B0(\key_mem[1][63] ), .B1(n3979), 
        .Y(n1930) );
  AO22X1 U2336 ( .A0(n3970), .A1(n1490), .B0(\key_mem[1][65] ), .B1(n3979), 
        .Y(n1928) );
  AO22X1 U2337 ( .A0(n3970), .A1(n1491), .B0(\key_mem[1][66] ), .B1(n3978), 
        .Y(n1927) );
  AO22X1 U2338 ( .A0(n3970), .A1(n1492), .B0(\key_mem[1][67] ), .B1(n3977), 
        .Y(n1926) );
  AO22X1 U2339 ( .A0(n3970), .A1(n1493), .B0(\key_mem[1][68] ), .B1(n3984), 
        .Y(n1925) );
  AO22X1 U2340 ( .A0(n3970), .A1(n1494), .B0(\key_mem[1][69] ), .B1(n3984), 
        .Y(n1924) );
  AO22X1 U2341 ( .A0(n3971), .A1(n1496), .B0(\key_mem[1][71] ), .B1(n3984), 
        .Y(n1922) );
  AO22X1 U2342 ( .A0(n3971), .A1(n1499), .B0(\key_mem[1][74] ), .B1(n3982), 
        .Y(n1919) );
  AO22X1 U2343 ( .A0(n3971), .A1(n1502), .B0(\key_mem[1][77] ), .B1(n3977), 
        .Y(n1916) );
  AO22X1 U2344 ( .A0(n3971), .A1(n1504), .B0(\key_mem[1][79] ), .B1(n3981), 
        .Y(n1914) );
  AO22X1 U2345 ( .A0(n3972), .A1(n1506), .B0(\key_mem[1][81] ), .B1(n3980), 
        .Y(n1912) );
  AO22X1 U2346 ( .A0(n3972), .A1(n1507), .B0(\key_mem[1][82] ), .B1(n3979), 
        .Y(n1911) );
  AO22X1 U2347 ( .A0(n3972), .A1(n1509), .B0(\key_mem[1][84] ), .B1(n3985), 
        .Y(n1909) );
  AO22X1 U2348 ( .A0(n3972), .A1(n1510), .B0(\key_mem[1][85] ), .B1(n3988), 
        .Y(n1908) );
  AO22X1 U2349 ( .A0(n3972), .A1(n1512), .B0(\key_mem[1][87] ), .B1(n3987), 
        .Y(n1906) );
  AO22X1 U2350 ( .A0(n3972), .A1(n1513), .B0(\key_mem[1][88] ), .B1(n3986), 
        .Y(n1905) );
  AO22X1 U2351 ( .A0(n3972), .A1(n1514), .B0(\key_mem[1][89] ), .B1(n3982), 
        .Y(n1904) );
  AO22X1 U2352 ( .A0(n3973), .A1(n1515), .B0(\key_mem[1][90] ), .B1(n3981), 
        .Y(n1903) );
  AO22X1 U2353 ( .A0(n3973), .A1(n1516), .B0(\key_mem[1][91] ), .B1(n3980), 
        .Y(n1902) );
  AO22X1 U2354 ( .A0(n3973), .A1(n1517), .B0(\key_mem[1][92] ), .B1(n3979), 
        .Y(n1901) );
  AO22X1 U2355 ( .A0(n3973), .A1(n1518), .B0(\key_mem[1][93] ), .B1(n3978), 
        .Y(n1900) );
  AO22X1 U2356 ( .A0(n3973), .A1(n1519), .B0(\key_mem[1][94] ), .B1(n3977), 
        .Y(n1899) );
  AO22X1 U2357 ( .A0(n3973), .A1(n1520), .B0(\key_mem[1][95] ), .B1(n3982), 
        .Y(n1898) );
  AO22X1 U2358 ( .A0(n3973), .A1(n1522), .B0(\key_mem[1][97] ), .B1(n3981), 
        .Y(n1896) );
  AO22X1 U2359 ( .A0(n3973), .A1(n1523), .B0(\key_mem[1][98] ), .B1(n3980), 
        .Y(n1895) );
  AO22X1 U2360 ( .A0(n3973), .A1(n1524), .B0(\key_mem[1][99] ), .B1(n3979), 
        .Y(n1894) );
  AO22X1 U2361 ( .A0(n3974), .A1(n1525), .B0(\key_mem[1][100] ), .B1(n3978), 
        .Y(n1893) );
  AO22X1 U2362 ( .A0(n3974), .A1(n1526), .B0(\key_mem[1][101] ), .B1(n3983), 
        .Y(n1892) );
  AO22X1 U2363 ( .A0(n3974), .A1(n1528), .B0(\key_mem[1][103] ), .B1(n3984), 
        .Y(n1890) );
  AO22X1 U2364 ( .A0(n3974), .A1(n1530), .B0(\key_mem[1][105] ), .B1(n3986), 
        .Y(n1888) );
  AO22X1 U2365 ( .A0(n3974), .A1(n1531), .B0(\key_mem[1][106] ), .B1(n3977), 
        .Y(n1887) );
  AO22X1 U2366 ( .A0(n3974), .A1(n1533), .B0(\key_mem[1][108] ), .B1(n3979), 
        .Y(n1885) );
  AO22X1 U2367 ( .A0(n3974), .A1(n1534), .B0(\key_mem[1][109] ), .B1(n3978), 
        .Y(n1884) );
  AO22X1 U2368 ( .A0(n3975), .A1(n1536), .B0(\key_mem[1][111] ), .B1(n3983), 
        .Y(n1882) );
  AO22X1 U2369 ( .A0(n3975), .A1(n1537), .B0(\key_mem[1][112] ), .B1(n3988), 
        .Y(n1881) );
  AO22X1 U2370 ( .A0(n3975), .A1(n1538), .B0(\key_mem[1][113] ), .B1(n3987), 
        .Y(n1880) );
  AO22X1 U2371 ( .A0(n3975), .A1(n1539), .B0(\key_mem[1][114] ), .B1(n3988), 
        .Y(n1879) );
  AO22X1 U2372 ( .A0(n3975), .A1(n1541), .B0(\key_mem[1][116] ), .B1(n3986), 
        .Y(n1877) );
  AO22X1 U2373 ( .A0(n3975), .A1(n1542), .B0(\key_mem[1][117] ), .B1(n3985), 
        .Y(n1876) );
  AO22X1 U2374 ( .A0(n3975), .A1(n1543), .B0(\key_mem[1][118] ), .B1(n3984), 
        .Y(n1875) );
  AO22X1 U2375 ( .A0(n3975), .A1(n1544), .B0(\key_mem[1][119] ), .B1(n3983), 
        .Y(n1874) );
  AO22X1 U2376 ( .A0(n3976), .A1(n1545), .B0(\key_mem[1][120] ), .B1(n3982), 
        .Y(n1873) );
  AO22X1 U2377 ( .A0(n3976), .A1(n1546), .B0(\key_mem[1][121] ), .B1(n3981), 
        .Y(n1872) );
  AO22X1 U2378 ( .A0(n3976), .A1(n1547), .B0(\key_mem[1][122] ), .B1(n3980), 
        .Y(n1871) );
  AO22X1 U2379 ( .A0(n3976), .A1(n1548), .B0(\key_mem[1][123] ), .B1(n3979), 
        .Y(n1870) );
  AO22X1 U2380 ( .A0(n3976), .A1(n1549), .B0(\key_mem[1][124] ), .B1(n3978), 
        .Y(n1869) );
  AO22X1 U2381 ( .A0(n3976), .A1(n1550), .B0(\key_mem[1][125] ), .B1(n3977), 
        .Y(n1868) );
  AO22X1 U2382 ( .A0(n3976), .A1(n1551), .B0(\key_mem[1][126] ), .B1(n3988), 
        .Y(n1867) );
  AO22X1 U2383 ( .A0(n3976), .A1(n1552), .B0(\key_mem[1][127] ), .B1(n3978), 
        .Y(n1866) );
  AO22X1 U2384 ( .A0(n4036), .A1(n1450), .B0(\key_mem[13][25] ), .B1(n4053), 
        .Y(n3504) );
  AO22X1 U2385 ( .A0(n4092), .A1(n695), .B0(\key_mem[11][25] ), .B1(n4107), 
        .Y(n3248) );
  AO22X1 U2386 ( .A0(n4148), .A1(n695), .B0(\key_mem[9][25] ), .B1(n4171), .Y(
        n2992) );
  AO22X1 U2387 ( .A0(n4205), .A1(n695), .B0(\key_mem[7][25] ), .B1(n4222), .Y(
        n2736) );
  AO22X1 U2388 ( .A0(n4260), .A1(n695), .B0(\key_mem[5][25] ), .B1(n4285), .Y(
        n2480) );
  AO22X1 U2389 ( .A0(n4316), .A1(n695), .B0(\key_mem[3][25] ), .B1(n4332), .Y(
        n2224) );
  AO22X1 U2390 ( .A0(n4039), .A1(n1482), .B0(\key_mem[13][57] ), .B1(n4053), 
        .Y(n3472) );
  AO22X1 U2391 ( .A0(n4095), .A1(n663), .B0(\key_mem[11][57] ), .B1(n4116), 
        .Y(n3216) );
  AO22X1 U2392 ( .A0(n4151), .A1(n663), .B0(\key_mem[9][57] ), .B1(n4166), .Y(
        n2960) );
  AO22X1 U2393 ( .A0(n4207), .A1(n663), .B0(\key_mem[7][57] ), .B1(n4220), .Y(
        n2704) );
  AO22X1 U2394 ( .A0(n4263), .A1(n663), .B0(\key_mem[5][57] ), .B1(n4285), .Y(
        n2448) );
  AO22X1 U2395 ( .A0(n4319), .A1(n663), .B0(\key_mem[3][57] ), .B1(n4340), .Y(
        n2192) );
  AO22X1 U2396 ( .A0(n4042), .A1(n1514), .B0(\key_mem[13][89] ), .B1(n4050), 
        .Y(n3440) );
  AO22X1 U2397 ( .A0(n4098), .A1(n631), .B0(\key_mem[11][89] ), .B1(n4105), 
        .Y(n3184) );
  AO22X1 U2398 ( .A0(n4154), .A1(n631), .B0(\key_mem[9][89] ), .B1(n4169), .Y(
        n2928) );
  AO22X1 U2399 ( .A0(n4210), .A1(n631), .B0(\key_mem[7][89] ), .B1(n4226), .Y(
        n2672) );
  AO22X1 U2400 ( .A0(n4266), .A1(n631), .B0(\key_mem[5][89] ), .B1(n4281), .Y(
        n2416) );
  AO22X1 U2401 ( .A0(n4322), .A1(n631), .B0(\key_mem[3][89] ), .B1(n4330), .Y(
        n2160) );
  AO22X1 U2402 ( .A0(n4046), .A1(n1546), .B0(\key_mem[13][121] ), .B1(n4053), 
        .Y(n3408) );
  AO22X1 U2403 ( .A0(n4102), .A1(n599), .B0(\key_mem[11][121] ), .B1(n4104), 
        .Y(n3152) );
  AO22X1 U2404 ( .A0(n4158), .A1(n599), .B0(\key_mem[9][121] ), .B1(n4167), 
        .Y(n2896) );
  AO22X1 U2405 ( .A0(n4202), .A1(n599), .B0(\key_mem[7][121] ), .B1(n4225), 
        .Y(n2640) );
  AO22X1 U2406 ( .A0(n4270), .A1(n599), .B0(\key_mem[5][121] ), .B1(n4279), 
        .Y(n2384) );
  AO22X1 U2407 ( .A0(n4326), .A1(n599), .B0(\key_mem[3][121] ), .B1(n4332), 
        .Y(n2128) );
  AO22X1 U2408 ( .A0(n4036), .A1(n1453), .B0(\key_mem[13][28] ), .B1(n4052), 
        .Y(n3501) );
  AO22X1 U2409 ( .A0(n4092), .A1(n692), .B0(\key_mem[11][28] ), .B1(n4116), 
        .Y(n3245) );
  AO22X1 U2410 ( .A0(n4148), .A1(n692), .B0(\key_mem[9][28] ), .B1(n4164), .Y(
        n2989) );
  AO22X1 U2411 ( .A0(n4205), .A1(n692), .B0(\key_mem[7][28] ), .B1(n4222), .Y(
        n2733) );
  AO22X1 U2412 ( .A0(n4260), .A1(n692), .B0(\key_mem[5][28] ), .B1(n4276), .Y(
        n2477) );
  AO22X1 U2413 ( .A0(n4316), .A1(n692), .B0(\key_mem[3][28] ), .B1(n4331), .Y(
        n2221) );
  AO22X1 U2414 ( .A0(n4040), .A1(n1485), .B0(\key_mem[13][60] ), .B1(n4052), 
        .Y(n3469) );
  AO22X1 U2415 ( .A0(n4096), .A1(n660), .B0(\key_mem[11][60] ), .B1(n4109), 
        .Y(n3213) );
  AO22X1 U2416 ( .A0(n4152), .A1(n660), .B0(\key_mem[9][60] ), .B1(n4165), .Y(
        n2957) );
  AO22X1 U2417 ( .A0(n4208), .A1(n660), .B0(\key_mem[7][60] ), .B1(n4228), .Y(
        n2701) );
  AO22X1 U2418 ( .A0(n4264), .A1(n660), .B0(\key_mem[5][60] ), .B1(n4281), .Y(
        n2445) );
  AO22X1 U2419 ( .A0(n4320), .A1(n660), .B0(\key_mem[3][60] ), .B1(n4328), .Y(
        n2189) );
  AO22X1 U2420 ( .A0(n4043), .A1(n1517), .B0(\key_mem[13][92] ), .B1(n4059), 
        .Y(n3437) );
  AO22X1 U2421 ( .A0(n4099), .A1(n628), .B0(\key_mem[11][92] ), .B1(n4107), 
        .Y(n3181) );
  AO22X1 U2422 ( .A0(n4155), .A1(n628), .B0(\key_mem[9][92] ), .B1(n4170), .Y(
        n2925) );
  AO22X1 U2423 ( .A0(n4211), .A1(n628), .B0(\key_mem[7][92] ), .B1(n4216), .Y(
        n2669) );
  AO22X1 U2424 ( .A0(n4267), .A1(n628), .B0(\key_mem[5][92] ), .B1(n4282), .Y(
        n2413) );
  AO22X1 U2425 ( .A0(n4323), .A1(n628), .B0(\key_mem[3][92] ), .B1(n4341), .Y(
        n2157) );
  AO22X1 U2426 ( .A0(n4046), .A1(n1549), .B0(\key_mem[13][124] ), .B1(n4052), 
        .Y(n3405) );
  AO22X1 U2427 ( .A0(n4102), .A1(n596), .B0(\key_mem[11][124] ), .B1(n4109), 
        .Y(n3149) );
  AO22X1 U2428 ( .A0(n4158), .A1(n596), .B0(\key_mem[9][124] ), .B1(n4167), 
        .Y(n2893) );
  AO22X1 U2429 ( .A0(n4202), .A1(n596), .B0(\key_mem[7][124] ), .B1(n4228), 
        .Y(n2637) );
  AO22X1 U2430 ( .A0(n4270), .A1(n596), .B0(\key_mem[5][124] ), .B1(n4279), 
        .Y(n2381) );
  AO22X1 U2431 ( .A0(n4326), .A1(n596), .B0(\key_mem[3][124] ), .B1(n4337), 
        .Y(n2125) );
  AO22X1 U2432 ( .A0(n4036), .A1(n1454), .B0(\key_mem[13][29] ), .B1(n4051), 
        .Y(n3500) );
  AO22X1 U2433 ( .A0(n4092), .A1(n691), .B0(\key_mem[11][29] ), .B1(n4105), 
        .Y(n3244) );
  AO22X1 U2434 ( .A0(n4148), .A1(n691), .B0(\key_mem[9][29] ), .B1(n4171), .Y(
        n2988) );
  AO22X1 U2435 ( .A0(n4205), .A1(n691), .B0(\key_mem[7][29] ), .B1(n4222), .Y(
        n2732) );
  AO22X1 U2436 ( .A0(n4260), .A1(n691), .B0(\key_mem[5][29] ), .B1(n4283), .Y(
        n2476) );
  AO22X1 U2437 ( .A0(n4316), .A1(n691), .B0(\key_mem[3][29] ), .B1(n4334), .Y(
        n2220) );
  AO22X1 U2438 ( .A0(n4040), .A1(n1486), .B0(\key_mem[13][61] ), .B1(n4055), 
        .Y(n3468) );
  AO22X1 U2439 ( .A0(n4096), .A1(n659), .B0(\key_mem[11][61] ), .B1(n4115), 
        .Y(n3212) );
  AO22X1 U2440 ( .A0(n4152), .A1(n659), .B0(\key_mem[9][61] ), .B1(n4170), .Y(
        n2956) );
  AO22X1 U2441 ( .A0(n4208), .A1(n659), .B0(\key_mem[7][61] ), .B1(n4227), .Y(
        n2700) );
  AO22X1 U2442 ( .A0(n4264), .A1(n659), .B0(\key_mem[5][61] ), .B1(n4273), .Y(
        n2444) );
  AO22X1 U2443 ( .A0(n4320), .A1(n659), .B0(\key_mem[3][61] ), .B1(n4332), .Y(
        n2188) );
  AO22X1 U2444 ( .A0(n4043), .A1(n1518), .B0(\key_mem[13][93] ), .B1(n4057), 
        .Y(n3436) );
  AO22X1 U2445 ( .A0(n4099), .A1(n627), .B0(\key_mem[11][93] ), .B1(n4106), 
        .Y(n3180) );
  AO22X1 U2446 ( .A0(n4155), .A1(n627), .B0(\key_mem[9][93] ), .B1(n4169), .Y(
        n2924) );
  AO22X1 U2447 ( .A0(n4211), .A1(n627), .B0(\key_mem[7][93] ), .B1(n4219), .Y(
        n2668) );
  AO22X1 U2448 ( .A0(n4267), .A1(n627), .B0(\key_mem[5][93] ), .B1(n4281), .Y(
        n2412) );
  AO22X1 U2449 ( .A0(n4323), .A1(n627), .B0(\key_mem[3][93] ), .B1(n4341), .Y(
        n2156) );
  AO22X1 U2450 ( .A0(n4046), .A1(n1550), .B0(\key_mem[13][125] ), .B1(n4051), 
        .Y(n3404) );
  AO22X1 U2451 ( .A0(n4102), .A1(n595), .B0(\key_mem[11][125] ), .B1(n4111), 
        .Y(n3148) );
  AO22X1 U2452 ( .A0(n4158), .A1(n595), .B0(\key_mem[9][125] ), .B1(n4166), 
        .Y(n2892) );
  AO22X1 U2453 ( .A0(n732), .A1(n595), .B0(\key_mem[7][125] ), .B1(n4228), .Y(
        n2636) );
  AO22X1 U2454 ( .A0(n4270), .A1(n595), .B0(\key_mem[5][125] ), .B1(n4278), 
        .Y(n2380) );
  AO22X1 U2455 ( .A0(n4326), .A1(n595), .B0(\key_mem[3][125] ), .B1(n4337), 
        .Y(n2124) );
  AO22X1 U2456 ( .A0(n4037), .A1(n1455), .B0(\key_mem[13][30] ), .B1(n4050), 
        .Y(n3499) );
  AO22X1 U2457 ( .A0(n4093), .A1(n690), .B0(\key_mem[11][30] ), .B1(n4116), 
        .Y(n3243) );
  AO22X1 U2458 ( .A0(n4149), .A1(n690), .B0(\key_mem[9][30] ), .B1(n4172), .Y(
        n2987) );
  AO22X1 U2459 ( .A0(n4206), .A1(n690), .B0(\key_mem[7][30] ), .B1(n4222), .Y(
        n2731) );
  AO22X1 U2460 ( .A0(n4261), .A1(n690), .B0(\key_mem[5][30] ), .B1(n4284), .Y(
        n2475) );
  AO22X1 U2461 ( .A0(n4317), .A1(n690), .B0(\key_mem[3][30] ), .B1(n4329), .Y(
        n2219) );
  AO22X1 U2462 ( .A0(n4040), .A1(n1487), .B0(\key_mem[13][62] ), .B1(n4059), 
        .Y(n3467) );
  AO22X1 U2463 ( .A0(n4096), .A1(n658), .B0(\key_mem[11][62] ), .B1(n4116), 
        .Y(n3211) );
  AO22X1 U2464 ( .A0(n4152), .A1(n658), .B0(\key_mem[9][62] ), .B1(n4169), .Y(
        n2955) );
  AO22X1 U2465 ( .A0(n4208), .A1(n658), .B0(\key_mem[7][62] ), .B1(n4227), .Y(
        n2699) );
  AO22X1 U2466 ( .A0(n4264), .A1(n658), .B0(\key_mem[5][62] ), .B1(n4272), .Y(
        n2443) );
  AO22X1 U2467 ( .A0(n4320), .A1(n658), .B0(\key_mem[3][62] ), .B1(n4338), .Y(
        n2187) );
  AO22X1 U2468 ( .A0(n4043), .A1(n1519), .B0(\key_mem[13][94] ), .B1(n4057), 
        .Y(n3435) );
  AO22X1 U2469 ( .A0(n4099), .A1(n626), .B0(\key_mem[11][94] ), .B1(n4113), 
        .Y(n3179) );
  AO22X1 U2470 ( .A0(n4155), .A1(n626), .B0(\key_mem[9][94] ), .B1(n4168), .Y(
        n2923) );
  AO22X1 U2471 ( .A0(n4211), .A1(n626), .B0(\key_mem[7][94] ), .B1(n4216), .Y(
        n2667) );
  AO22X1 U2472 ( .A0(n4267), .A1(n626), .B0(\key_mem[5][94] ), .B1(n4280), .Y(
        n2411) );
  AO22X1 U2473 ( .A0(n4323), .A1(n626), .B0(\key_mem[3][94] ), .B1(n4339), .Y(
        n2155) );
  AO22X1 U2474 ( .A0(n4046), .A1(n1551), .B0(\key_mem[13][126] ), .B1(n4050), 
        .Y(n3403) );
  AO22X1 U2475 ( .A0(n4102), .A1(n594), .B0(\key_mem[11][126] ), .B1(n4108), 
        .Y(n3147) );
  AO22X1 U2476 ( .A0(n4158), .A1(n594), .B0(\key_mem[9][126] ), .B1(n4165), 
        .Y(n2891) );
  AO22X1 U2477 ( .A0(n732), .A1(n594), .B0(\key_mem[7][126] ), .B1(n4229), .Y(
        n2635) );
  AO22X1 U2478 ( .A0(n4270), .A1(n594), .B0(\key_mem[5][126] ), .B1(n4277), 
        .Y(n2379) );
  AO22X1 U2479 ( .A0(n4326), .A1(n594), .B0(\key_mem[3][126] ), .B1(n4337), 
        .Y(n2123) );
  AO22X1 U2480 ( .A0(n4036), .A1(n1452), .B0(\key_mem[13][27] ), .B1(n4058), 
        .Y(n3502) );
  AO22X1 U2481 ( .A0(n4092), .A1(n693), .B0(\key_mem[11][27] ), .B1(n4117), 
        .Y(n3246) );
  AO22X1 U2482 ( .A0(n4148), .A1(n693), .B0(\key_mem[9][27] ), .B1(n4173), .Y(
        n2990) );
  AO22X1 U2483 ( .A0(n4205), .A1(n693), .B0(\key_mem[7][27] ), .B1(n4222), .Y(
        n2734) );
  AO22X1 U2484 ( .A0(n4260), .A1(n693), .B0(\key_mem[5][27] ), .B1(n4285), .Y(
        n2478) );
  AO22X1 U2485 ( .A0(n4316), .A1(n693), .B0(\key_mem[3][27] ), .B1(n4328), .Y(
        n2222) );
  AO22X1 U2486 ( .A0(n4039), .A1(n1484), .B0(\key_mem[13][59] ), .B1(n4060), 
        .Y(n3470) );
  AO22X1 U2487 ( .A0(n4095), .A1(n661), .B0(\key_mem[11][59] ), .B1(n4117), 
        .Y(n3214) );
  AO22X1 U2488 ( .A0(n4151), .A1(n661), .B0(\key_mem[9][59] ), .B1(n4161), .Y(
        n2958) );
  AO22X1 U2489 ( .A0(n4207), .A1(n661), .B0(\key_mem[7][59] ), .B1(n4217), .Y(
        n2702) );
  AO22X1 U2490 ( .A0(n4263), .A1(n661), .B0(\key_mem[5][59] ), .B1(n4277), .Y(
        n2446) );
  AO22X1 U2491 ( .A0(n4319), .A1(n661), .B0(\key_mem[3][59] ), .B1(n4340), .Y(
        n2190) );
  AO22X1 U2492 ( .A0(n4043), .A1(n1516), .B0(\key_mem[13][91] ), .B1(n4050), 
        .Y(n3438) );
  AO22X1 U2493 ( .A0(n4099), .A1(n629), .B0(\key_mem[11][91] ), .B1(n4105), 
        .Y(n3182) );
  AO22X1 U2494 ( .A0(n4155), .A1(n629), .B0(\key_mem[9][91] ), .B1(n4169), .Y(
        n2926) );
  AO22X1 U2495 ( .A0(n4211), .A1(n629), .B0(\key_mem[7][91] ), .B1(n4217), .Y(
        n2670) );
  AO22X1 U2496 ( .A0(n4267), .A1(n629), .B0(\key_mem[5][91] ), .B1(n4281), .Y(
        n2414) );
  AO22X1 U2497 ( .A0(n4323), .A1(n629), .B0(\key_mem[3][91] ), .B1(n4339), .Y(
        n2158) );
  AO22X1 U2498 ( .A0(n4046), .A1(n1548), .B0(\key_mem[13][123] ), .B1(n4049), 
        .Y(n3406) );
  AO22X1 U2499 ( .A0(n4102), .A1(n597), .B0(\key_mem[11][123] ), .B1(n4104), 
        .Y(n3150) );
  AO22X1 U2500 ( .A0(n4158), .A1(n597), .B0(\key_mem[9][123] ), .B1(n4161), 
        .Y(n2894) );
  AO22X1 U2501 ( .A0(n732), .A1(n597), .B0(\key_mem[7][123] ), .B1(n4226), .Y(
        n2638) );
  AO22X1 U2502 ( .A0(n4270), .A1(n597), .B0(\key_mem[5][123] ), .B1(n4273), 
        .Y(n2382) );
  AO22X1 U2503 ( .A0(n4326), .A1(n597), .B0(\key_mem[3][123] ), .B1(n4337), 
        .Y(n2126) );
  AO22X1 U2504 ( .A0(n4036), .A1(n1451), .B0(\key_mem[13][26] ), .B1(n4054), 
        .Y(n3503) );
  AO22X1 U2505 ( .A0(n4092), .A1(n694), .B0(\key_mem[11][26] ), .B1(n4111), 
        .Y(n3247) );
  AO22X1 U2506 ( .A0(n4148), .A1(n694), .B0(\key_mem[9][26] ), .B1(n4172), .Y(
        n2991) );
  AO22X1 U2507 ( .A0(n4205), .A1(n694), .B0(\key_mem[7][26] ), .B1(n4222), .Y(
        n2735) );
  AO22X1 U2508 ( .A0(n4260), .A1(n694), .B0(\key_mem[5][26] ), .B1(n4284), .Y(
        n2479) );
  AO22X1 U2509 ( .A0(n4316), .A1(n694), .B0(\key_mem[3][26] ), .B1(n4331), .Y(
        n2223) );
  AO22X1 U2510 ( .A0(n4039), .A1(n1483), .B0(\key_mem[13][58] ), .B1(n4061), 
        .Y(n3471) );
  AO22X1 U2511 ( .A0(n4095), .A1(n662), .B0(\key_mem[11][58] ), .B1(n4105), 
        .Y(n3215) );
  AO22X1 U2512 ( .A0(n4151), .A1(n662), .B0(\key_mem[9][58] ), .B1(n4159), .Y(
        n2959) );
  AO22X1 U2513 ( .A0(n4207), .A1(n662), .B0(\key_mem[7][58] ), .B1(n4215), .Y(
        n2703) );
  AO22X1 U2514 ( .A0(n4263), .A1(n662), .B0(\key_mem[5][58] ), .B1(n4271), .Y(
        n2447) );
  AO22X1 U2515 ( .A0(n4319), .A1(n662), .B0(\key_mem[3][58] ), .B1(n4330), .Y(
        n2191) );
  AO22X1 U2516 ( .A0(n4043), .A1(n1515), .B0(\key_mem[13][90] ), .B1(n4061), 
        .Y(n3439) );
  AO22X1 U2517 ( .A0(n4099), .A1(n630), .B0(\key_mem[11][90] ), .B1(n4107), 
        .Y(n3183) );
  AO22X1 U2518 ( .A0(n4155), .A1(n630), .B0(\key_mem[9][90] ), .B1(n4168), .Y(
        n2927) );
  AO22X1 U2519 ( .A0(n4211), .A1(n630), .B0(\key_mem[7][90] ), .B1(n4214), .Y(
        n2671) );
  AO22X1 U2520 ( .A0(n4267), .A1(n630), .B0(\key_mem[5][90] ), .B1(n4280), .Y(
        n2415) );
  AO22X1 U2521 ( .A0(n4323), .A1(n630), .B0(\key_mem[3][90] ), .B1(n4340), .Y(
        n2159) );
  AO22X1 U2522 ( .A0(n4046), .A1(n1547), .B0(\key_mem[13][122] ), .B1(n4052), 
        .Y(n3407) );
  AO22X1 U2523 ( .A0(n4102), .A1(n598), .B0(\key_mem[11][122] ), .B1(n4117), 
        .Y(n3151) );
  AO22X1 U2524 ( .A0(n4158), .A1(n598), .B0(\key_mem[9][122] ), .B1(n4166), 
        .Y(n2895) );
  AO22X1 U2525 ( .A0(n732), .A1(n598), .B0(\key_mem[7][122] ), .B1(n4225), .Y(
        n2639) );
  AO22X1 U2526 ( .A0(n4270), .A1(n598), .B0(\key_mem[5][122] ), .B1(n4278), 
        .Y(n2383) );
  AO22X1 U2527 ( .A0(n4326), .A1(n598), .B0(\key_mem[3][122] ), .B1(n4333), 
        .Y(n2127) );
  AO22X1 U2528 ( .A0(n4036), .A1(n1449), .B0(\key_mem[13][24] ), .B1(n4053), 
        .Y(n3505) );
  AO22X1 U2529 ( .A0(n4092), .A1(n696), .B0(\key_mem[11][24] ), .B1(n4109), 
        .Y(n3249) );
  AO22X1 U2530 ( .A0(n4148), .A1(n696), .B0(\key_mem[9][24] ), .B1(n4162), .Y(
        n2993) );
  AO22X1 U2531 ( .A0(n4205), .A1(n696), .B0(\key_mem[7][24] ), .B1(n4222), .Y(
        n2737) );
  AO22X1 U2532 ( .A0(n4260), .A1(n696), .B0(\key_mem[5][24] ), .B1(n4274), .Y(
        n2481) );
  AO22X1 U2533 ( .A0(n4316), .A1(n696), .B0(\key_mem[3][24] ), .B1(n4327), .Y(
        n2225) );
  AO22X1 U2534 ( .A0(n4039), .A1(n1481), .B0(\key_mem[13][56] ), .B1(n4051), 
        .Y(n3473) );
  AO22X1 U2535 ( .A0(n4095), .A1(n664), .B0(\key_mem[11][56] ), .B1(n4106), 
        .Y(n3217) );
  AO22X1 U2536 ( .A0(n4151), .A1(n664), .B0(\key_mem[9][56] ), .B1(n4169), .Y(
        n2961) );
  AO22X1 U2537 ( .A0(n4207), .A1(n664), .B0(\key_mem[7][56] ), .B1(n4217), .Y(
        n2705) );
  AO22X1 U2538 ( .A0(n4263), .A1(n664), .B0(\key_mem[5][56] ), .B1(n4281), .Y(
        n2449) );
  AO22X1 U2539 ( .A0(n4319), .A1(n664), .B0(\key_mem[3][56] ), .B1(n4328), .Y(
        n2193) );
  AO22X1 U2540 ( .A0(n4042), .A1(n1513), .B0(\key_mem[13][88] ), .B1(n4060), 
        .Y(n3441) );
  AO22X1 U2541 ( .A0(n4098), .A1(n632), .B0(\key_mem[11][88] ), .B1(n4112), 
        .Y(n3185) );
  AO22X1 U2542 ( .A0(n4154), .A1(n632), .B0(\key_mem[9][88] ), .B1(n4159), .Y(
        n2929) );
  AO22X1 U2543 ( .A0(n4210), .A1(n632), .B0(\key_mem[7][88] ), .B1(n4215), .Y(
        n2673) );
  AO22X1 U2544 ( .A0(n4266), .A1(n632), .B0(\key_mem[5][88] ), .B1(n4278), .Y(
        n2417) );
  AO22X1 U2545 ( .A0(n4322), .A1(n632), .B0(\key_mem[3][88] ), .B1(n725), .Y(
        n2161) );
  AO22X1 U2546 ( .A0(n4046), .A1(n1545), .B0(\key_mem[13][120] ), .B1(n4051), 
        .Y(n3409) );
  AO22X1 U2547 ( .A0(n4102), .A1(n600), .B0(\key_mem[11][120] ), .B1(n4108), 
        .Y(n3153) );
  AO22X1 U2548 ( .A0(n4158), .A1(n600), .B0(\key_mem[9][120] ), .B1(n4165), 
        .Y(n2897) );
  AO22X1 U2549 ( .A0(n732), .A1(n600), .B0(\key_mem[7][120] ), .B1(n4225), .Y(
        n2641) );
  AO22X1 U2550 ( .A0(n4270), .A1(n600), .B0(\key_mem[5][120] ), .B1(n4277), 
        .Y(n2385) );
  AO22X1 U2551 ( .A0(n4326), .A1(n600), .B0(\key_mem[3][120] ), .B1(n4331), 
        .Y(n2129) );
  AO22X1 U2552 ( .A0(n4037), .A1(n1456), .B0(\key_mem[13][31] ), .B1(n4052), 
        .Y(n3498) );
  AO22X1 U2553 ( .A0(n4093), .A1(n689), .B0(\key_mem[11][31] ), .B1(n4105), 
        .Y(n3242) );
  AO22X1 U2554 ( .A0(n4149), .A1(n689), .B0(\key_mem[9][31] ), .B1(n4167), .Y(
        n2986) );
  AO22X1 U2555 ( .A0(n4206), .A1(n689), .B0(\key_mem[7][31] ), .B1(n4222), .Y(
        n2730) );
  AO22X1 U2556 ( .A0(n4261), .A1(n689), .B0(\key_mem[5][31] ), .B1(n4283), .Y(
        n2474) );
  AO22X1 U2557 ( .A0(n4317), .A1(n689), .B0(\key_mem[3][31] ), .B1(n4335), .Y(
        n2218) );
  AO22X1 U2558 ( .A0(n4040), .A1(n1488), .B0(\key_mem[13][63] ), .B1(n4058), 
        .Y(n3466) );
  AO22X1 U2559 ( .A0(n4096), .A1(n657), .B0(\key_mem[11][63] ), .B1(n4109), 
        .Y(n3210) );
  AO22X1 U2560 ( .A0(n4152), .A1(n657), .B0(\key_mem[9][63] ), .B1(n4167), .Y(
        n2954) );
  AO22X1 U2561 ( .A0(n4208), .A1(n657), .B0(\key_mem[7][63] ), .B1(n4214), .Y(
        n2698) );
  AO22X1 U2562 ( .A0(n4264), .A1(n657), .B0(\key_mem[5][63] ), .B1(n4277), .Y(
        n2442) );
  AO22X1 U2563 ( .A0(n4320), .A1(n657), .B0(\key_mem[3][63] ), .B1(n4335), .Y(
        n2186) );
  AO22X1 U2564 ( .A0(n4043), .A1(n1520), .B0(\key_mem[13][95] ), .B1(n4057), 
        .Y(n3434) );
  AO22X1 U2565 ( .A0(n4099), .A1(n625), .B0(\key_mem[11][95] ), .B1(n4112), 
        .Y(n3178) );
  AO22X1 U2566 ( .A0(n4155), .A1(n625), .B0(\key_mem[9][95] ), .B1(n4170), .Y(
        n2922) );
  AO22X1 U2567 ( .A0(n4211), .A1(n625), .B0(\key_mem[7][95] ), .B1(n4218), .Y(
        n2666) );
  AO22X1 U2568 ( .A0(n4267), .A1(n625), .B0(\key_mem[5][95] ), .B1(n4282), .Y(
        n2410) );
  AO22X1 U2569 ( .A0(n4323), .A1(n625), .B0(\key_mem[3][95] ), .B1(n4340), .Y(
        n2154) );
  AO22X1 U2570 ( .A0(n4046), .A1(n1552), .B0(\key_mem[13][127] ), .B1(n4054), 
        .Y(n3402) );
  AO22X1 U2571 ( .A0(n4102), .A1(n593), .B0(\key_mem[11][127] ), .B1(n4106), 
        .Y(n3146) );
  AO22X1 U2572 ( .A0(n4158), .A1(n593), .B0(\key_mem[9][127] ), .B1(n4170), 
        .Y(n2890) );
  AO22X1 U2573 ( .A0(n732), .A1(n593), .B0(\key_mem[7][127] ), .B1(n4226), .Y(
        n2634) );
  AO22X1 U2574 ( .A0(n4270), .A1(n593), .B0(\key_mem[5][127] ), .B1(n4282), 
        .Y(n2378) );
  AO22X1 U2575 ( .A0(n4326), .A1(n593), .B0(\key_mem[3][127] ), .B1(n4337), 
        .Y(n2122) );
  AO22X1 U2576 ( .A0(n4034), .A1(n1426), .B0(\key_mem[13][1] ), .B1(n4047), 
        .Y(n3528) );
  AO22X1 U2577 ( .A0(n4090), .A1(n719), .B0(\key_mem[11][1] ), .B1(n4103), .Y(
        n3272) );
  AO22X1 U2578 ( .A0(n4146), .A1(n719), .B0(\key_mem[9][1] ), .B1(n4159), .Y(
        n3016) );
  AO22X1 U2579 ( .A0(n4203), .A1(n719), .B0(\key_mem[7][1] ), .B1(n4214), .Y(
        n2760) );
  AO22X1 U2580 ( .A0(n4258), .A1(n719), .B0(\key_mem[5][1] ), .B1(n4271), .Y(
        n2504) );
  AO22X1 U2581 ( .A0(n4314), .A1(n719), .B0(\key_mem[3][1] ), .B1(n4327), .Y(
        n2248) );
  AO22X1 U2582 ( .A0(n4034), .A1(n1427), .B0(\key_mem[13][2] ), .B1(n4048), 
        .Y(n3527) );
  AO22X1 U2583 ( .A0(n4090), .A1(n718), .B0(\key_mem[11][2] ), .B1(n4104), .Y(
        n3271) );
  AO22X1 U2584 ( .A0(n4146), .A1(n718), .B0(\key_mem[9][2] ), .B1(n4160), .Y(
        n3015) );
  AO22X1 U2585 ( .A0(n4203), .A1(n718), .B0(\key_mem[7][2] ), .B1(n4227), .Y(
        n2759) );
  AO22X1 U2586 ( .A0(n4258), .A1(n718), .B0(\key_mem[5][2] ), .B1(n4272), .Y(
        n2503) );
  AO22X1 U2587 ( .A0(n4314), .A1(n718), .B0(\key_mem[3][2] ), .B1(n4328), .Y(
        n2247) );
  AO22X1 U2588 ( .A0(n4034), .A1(n1428), .B0(\key_mem[13][3] ), .B1(n4049), 
        .Y(n3526) );
  AO22X1 U2589 ( .A0(n4090), .A1(n717), .B0(\key_mem[11][3] ), .B1(n4105), .Y(
        n3270) );
  AO22X1 U2590 ( .A0(n4146), .A1(n717), .B0(\key_mem[9][3] ), .B1(n4161), .Y(
        n3014) );
  AO22X1 U2591 ( .A0(n4203), .A1(n717), .B0(\key_mem[7][3] ), .B1(n4228), .Y(
        n2758) );
  AO22X1 U2592 ( .A0(n4258), .A1(n717), .B0(\key_mem[5][3] ), .B1(n4273), .Y(
        n2502) );
  AO22X1 U2593 ( .A0(n4314), .A1(n717), .B0(\key_mem[3][3] ), .B1(n4329), .Y(
        n2246) );
  AO22X1 U2594 ( .A0(n4034), .A1(n1429), .B0(\key_mem[13][4] ), .B1(n4050), 
        .Y(n3525) );
  AO22X1 U2595 ( .A0(n4090), .A1(n1429), .B0(\key_mem[11][4] ), .B1(n4106), 
        .Y(n3269) );
  AO22X1 U2596 ( .A0(n4146), .A1(n1429), .B0(\key_mem[9][4] ), .B1(n4162), .Y(
        n3013) );
  AO22X1 U2597 ( .A0(n4203), .A1(n1429), .B0(\key_mem[7][4] ), .B1(n4214), .Y(
        n2757) );
  AO22X1 U2598 ( .A0(n4258), .A1(n1429), .B0(\key_mem[5][4] ), .B1(n4274), .Y(
        n2501) );
  AO22X1 U2599 ( .A0(n4314), .A1(n1429), .B0(\key_mem[3][4] ), .B1(n4330), .Y(
        n2245) );
  AO22X1 U2600 ( .A0(n4034), .A1(n1430), .B0(\key_mem[13][5] ), .B1(n4051), 
        .Y(n3524) );
  AO22X1 U2601 ( .A0(n4090), .A1(n715), .B0(\key_mem[11][5] ), .B1(n4107), .Y(
        n3268) );
  AO22X1 U2602 ( .A0(n4146), .A1(n715), .B0(\key_mem[9][5] ), .B1(n4163), .Y(
        n3012) );
  AO22X1 U2603 ( .A0(n4203), .A1(n715), .B0(\key_mem[7][5] ), .B1(n4214), .Y(
        n2756) );
  AO22X1 U2604 ( .A0(n4258), .A1(n715), .B0(\key_mem[5][5] ), .B1(n4275), .Y(
        n2500) );
  AO22X1 U2605 ( .A0(n4314), .A1(n715), .B0(\key_mem[3][5] ), .B1(n4331), .Y(
        n2244) );
  AO22X1 U2606 ( .A0(n4034), .A1(n1432), .B0(\key_mem[13][7] ), .B1(n4053), 
        .Y(n3522) );
  AO22X1 U2607 ( .A0(n4090), .A1(n713), .B0(\key_mem[11][7] ), .B1(n4109), .Y(
        n3266) );
  AO22X1 U2608 ( .A0(n4146), .A1(n713), .B0(\key_mem[9][7] ), .B1(n4165), .Y(
        n3010) );
  AO22X1 U2609 ( .A0(n4203), .A1(n713), .B0(\key_mem[7][7] ), .B1(n4215), .Y(
        n2754) );
  AO22X1 U2610 ( .A0(n4258), .A1(n713), .B0(\key_mem[5][7] ), .B1(n4277), .Y(
        n2498) );
  AO22X1 U2611 ( .A0(n4314), .A1(n713), .B0(\key_mem[3][7] ), .B1(n4333), .Y(
        n2242) );
  AO22X1 U2612 ( .A0(n4035), .A1(n1435), .B0(\key_mem[13][10] ), .B1(n4056), 
        .Y(n3519) );
  AO22X1 U2613 ( .A0(n4091), .A1(n710), .B0(\key_mem[11][10] ), .B1(n4112), 
        .Y(n3263) );
  AO22X1 U2614 ( .A0(n4147), .A1(n710), .B0(\key_mem[9][10] ), .B1(n4168), .Y(
        n3007) );
  AO22X1 U2615 ( .A0(n4204), .A1(n710), .B0(\key_mem[7][10] ), .B1(n4218), .Y(
        n2751) );
  AO22X1 U2616 ( .A0(n4259), .A1(n710), .B0(\key_mem[5][10] ), .B1(n4280), .Y(
        n2495) );
  AO22X1 U2617 ( .A0(n4315), .A1(n710), .B0(\key_mem[3][10] ), .B1(n4330), .Y(
        n2239) );
  AO22X1 U2618 ( .A0(n4035), .A1(n1438), .B0(\key_mem[13][13] ), .B1(n4047), 
        .Y(n3516) );
  AO22X1 U2619 ( .A0(n4091), .A1(n707), .B0(\key_mem[11][13] ), .B1(n4103), 
        .Y(n3260) );
  AO22X1 U2620 ( .A0(n4147), .A1(n707), .B0(\key_mem[9][13] ), .B1(n4172), .Y(
        n3004) );
  AO22X1 U2621 ( .A0(n4204), .A1(n707), .B0(\key_mem[7][13] ), .B1(n4221), .Y(
        n2748) );
  AO22X1 U2622 ( .A0(n4259), .A1(n707), .B0(\key_mem[5][13] ), .B1(n4284), .Y(
        n2492) );
  AO22X1 U2623 ( .A0(n4315), .A1(n707), .B0(\key_mem[3][13] ), .B1(n4330), .Y(
        n2236) );
  AO22X1 U2624 ( .A0(n4035), .A1(n1443), .B0(\key_mem[13][18] ), .B1(n4048), 
        .Y(n3511) );
  AO22X1 U2625 ( .A0(n4091), .A1(n702), .B0(\key_mem[11][18] ), .B1(n4116), 
        .Y(n3255) );
  AO22X1 U2626 ( .A0(n4147), .A1(n702), .B0(\key_mem[9][18] ), .B1(n4173), .Y(
        n2999) );
  AO22X1 U2627 ( .A0(n4204), .A1(n702), .B0(\key_mem[7][18] ), .B1(n4221), .Y(
        n2743) );
  AO22X1 U2628 ( .A0(n4259), .A1(n702), .B0(\key_mem[5][18] ), .B1(n4285), .Y(
        n2487) );
  AO22X1 U2629 ( .A0(n4315), .A1(n702), .B0(\key_mem[3][18] ), .B1(n4339), .Y(
        n2231) );
  AO22X1 U2630 ( .A0(n4036), .A1(n1447), .B0(\key_mem[13][22] ), .B1(n4047), 
        .Y(n3507) );
  AO22X1 U2631 ( .A0(n4092), .A1(n698), .B0(\key_mem[11][22] ), .B1(n4117), 
        .Y(n3251) );
  AO22X1 U2632 ( .A0(n4148), .A1(n698), .B0(\key_mem[9][22] ), .B1(n4164), .Y(
        n2995) );
  AO22X1 U2633 ( .A0(n4205), .A1(n698), .B0(\key_mem[7][22] ), .B1(n4221), .Y(
        n2739) );
  AO22X1 U2634 ( .A0(n4260), .A1(n698), .B0(\key_mem[5][22] ), .B1(n4276), .Y(
        n2483) );
  AO22X1 U2635 ( .A0(n4316), .A1(n698), .B0(\key_mem[3][22] ), .B1(n4337), .Y(
        n2227) );
  AO22X1 U2636 ( .A0(n4037), .A1(n1458), .B0(\key_mem[13][33] ), .B1(n4060), 
        .Y(n3496) );
  AO22X1 U2637 ( .A0(n4093), .A1(n687), .B0(\key_mem[11][33] ), .B1(n4110), 
        .Y(n3240) );
  AO22X1 U2638 ( .A0(n4149), .A1(n687), .B0(\key_mem[9][33] ), .B1(n4163), .Y(
        n2984) );
  AO22X1 U2639 ( .A0(n4206), .A1(n687), .B0(\key_mem[7][33] ), .B1(n4223), .Y(
        n2728) );
  AO22X1 U2640 ( .A0(n4261), .A1(n687), .B0(\key_mem[5][33] ), .B1(n4274), .Y(
        n2472) );
  AO22X1 U2641 ( .A0(n4317), .A1(n687), .B0(\key_mem[3][33] ), .B1(n4330), .Y(
        n2216) );
  AO22X1 U2642 ( .A0(n4037), .A1(n1459), .B0(\key_mem[13][34] ), .B1(n4048), 
        .Y(n3495) );
  AO22X1 U2643 ( .A0(n4093), .A1(n686), .B0(\key_mem[11][34] ), .B1(n4115), 
        .Y(n3239) );
  AO22X1 U2644 ( .A0(n4149), .A1(n686), .B0(\key_mem[9][34] ), .B1(n4171), .Y(
        n2983) );
  AO22X1 U2645 ( .A0(n4206), .A1(n686), .B0(\key_mem[7][34] ), .B1(n4223), .Y(
        n2727) );
  AO22X1 U2646 ( .A0(n4261), .A1(n686), .B0(\key_mem[5][34] ), .B1(n4283), .Y(
        n2471) );
  AO22X1 U2647 ( .A0(n4317), .A1(n686), .B0(\key_mem[3][34] ), .B1(n4329), .Y(
        n2215) );
  AO22X1 U2648 ( .A0(n4037), .A1(n1460), .B0(\key_mem[13][35] ), .B1(n4053), 
        .Y(n3494) );
  AO22X1 U2649 ( .A0(n4093), .A1(n685), .B0(\key_mem[11][35] ), .B1(n4103), 
        .Y(n3238) );
  AO22X1 U2650 ( .A0(n4149), .A1(n685), .B0(\key_mem[9][35] ), .B1(n4172), .Y(
        n2982) );
  AO22X1 U2651 ( .A0(n4206), .A1(n685), .B0(\key_mem[7][35] ), .B1(n4223), .Y(
        n2726) );
  AO22X1 U2652 ( .A0(n4261), .A1(n685), .B0(\key_mem[5][35] ), .B1(n4284), .Y(
        n2470) );
  AO22X1 U2653 ( .A0(n4317), .A1(n685), .B0(\key_mem[3][35] ), .B1(n4333), .Y(
        n2214) );
  AO22X1 U2654 ( .A0(n4037), .A1(n1461), .B0(\key_mem[13][36] ), .B1(n4058), 
        .Y(n3493) );
  AO22X1 U2655 ( .A0(n4093), .A1(n684), .B0(\key_mem[11][36] ), .B1(n4116), 
        .Y(n3237) );
  AO22X1 U2656 ( .A0(n4149), .A1(n684), .B0(\key_mem[9][36] ), .B1(n4173), .Y(
        n2981) );
  AO22X1 U2657 ( .A0(n4206), .A1(n684), .B0(\key_mem[7][36] ), .B1(n4223), .Y(
        n2725) );
  AO22X1 U2658 ( .A0(n4261), .A1(n684), .B0(\key_mem[5][36] ), .B1(n4285), .Y(
        n2469) );
  AO22X1 U2659 ( .A0(n4317), .A1(n684), .B0(\key_mem[3][36] ), .B1(n4331), .Y(
        n2213) );
  AO22X1 U2660 ( .A0(n4037), .A1(n1462), .B0(\key_mem[13][37] ), .B1(n4059), 
        .Y(n3492) );
  AO22X1 U2661 ( .A0(n4093), .A1(n683), .B0(\key_mem[11][37] ), .B1(n4117), 
        .Y(n3236) );
  AO22X1 U2662 ( .A0(n4149), .A1(n683), .B0(\key_mem[9][37] ), .B1(n4172), .Y(
        n2980) );
  AO22X1 U2663 ( .A0(n4206), .A1(n683), .B0(\key_mem[7][37] ), .B1(n4223), .Y(
        n2724) );
  AO22X1 U2664 ( .A0(n4261), .A1(n683), .B0(\key_mem[5][37] ), .B1(n4283), .Y(
        n2468) );
  AO22X1 U2665 ( .A0(n4317), .A1(n683), .B0(\key_mem[3][37] ), .B1(n4327), .Y(
        n2212) );
  AO22X1 U2666 ( .A0(n4037), .A1(n1464), .B0(\key_mem[13][39] ), .B1(n4060), 
        .Y(n3490) );
  AO22X1 U2667 ( .A0(n4093), .A1(n681), .B0(\key_mem[11][39] ), .B1(n4109), 
        .Y(n3234) );
  AO22X1 U2668 ( .A0(n4149), .A1(n681), .B0(\key_mem[9][39] ), .B1(n4173), .Y(
        n2978) );
  AO22X1 U2669 ( .A0(n4206), .A1(n681), .B0(\key_mem[7][39] ), .B1(n4223), .Y(
        n2722) );
  AO22X1 U2670 ( .A0(n4261), .A1(n681), .B0(\key_mem[5][39] ), .B1(n4285), .Y(
        n2466) );
  AO22X1 U2671 ( .A0(n4317), .A1(n681), .B0(\key_mem[3][39] ), .B1(n4328), .Y(
        n2210) );
  AO22X1 U2672 ( .A0(n4038), .A1(n1467), .B0(\key_mem[13][42] ), .B1(n4054), 
        .Y(n3487) );
  AO22X1 U2673 ( .A0(n4094), .A1(n678), .B0(\key_mem[11][42] ), .B1(n4110), 
        .Y(n3231) );
  AO22X1 U2674 ( .A0(n4150), .A1(n678), .B0(\key_mem[9][42] ), .B1(n4166), .Y(
        n2975) );
  AO22X1 U2675 ( .A0(n732), .A1(n678), .B0(\key_mem[7][42] ), .B1(n4223), .Y(
        n2719) );
  AO22X1 U2676 ( .A0(n4262), .A1(n678), .B0(\key_mem[5][42] ), .B1(n4277), .Y(
        n2463) );
  AO22X1 U2677 ( .A0(n4318), .A1(n678), .B0(\key_mem[3][42] ), .B1(n4331), .Y(
        n2207) );
  AO22X1 U2678 ( .A0(n4038), .A1(n1470), .B0(\key_mem[13][45] ), .B1(n4059), 
        .Y(n3484) );
  AO22X1 U2679 ( .A0(n4094), .A1(n675), .B0(\key_mem[11][45] ), .B1(n4108), 
        .Y(n3228) );
  AO22X1 U2680 ( .A0(n4150), .A1(n675), .B0(\key_mem[9][45] ), .B1(n4159), .Y(
        n2972) );
  AO22X1 U2681 ( .A0(n4202), .A1(n675), .B0(\key_mem[7][45] ), .B1(n4214), .Y(
        n2716) );
  AO22X1 U2682 ( .A0(n4262), .A1(n675), .B0(\key_mem[5][45] ), .B1(n4272), .Y(
        n2460) );
  AO22X1 U2683 ( .A0(n4318), .A1(n675), .B0(\key_mem[3][45] ), .B1(n4341), .Y(
        n2204) );
  AO22X1 U2684 ( .A0(n4039), .A1(n1475), .B0(\key_mem[13][50] ), .B1(n4060), 
        .Y(n3479) );
  AO22X1 U2685 ( .A0(n4095), .A1(n670), .B0(\key_mem[11][50] ), .B1(n4110), 
        .Y(n3223) );
  AO22X1 U2686 ( .A0(n4151), .A1(n670), .B0(\key_mem[9][50] ), .B1(n4165), .Y(
        n2967) );
  AO22X1 U2687 ( .A0(n4207), .A1(n670), .B0(\key_mem[7][50] ), .B1(n4215), .Y(
        n2711) );
  AO22X1 U2688 ( .A0(n4263), .A1(n670), .B0(\key_mem[5][50] ), .B1(n4277), .Y(
        n2455) );
  AO22X1 U2689 ( .A0(n4319), .A1(n670), .B0(\key_mem[3][50] ), .B1(n4339), .Y(
        n2199) );
  AO22X1 U2690 ( .A0(n4039), .A1(n1478), .B0(\key_mem[13][53] ), .B1(n4049), 
        .Y(n3476) );
  AO22X1 U2691 ( .A0(n4095), .A1(n667), .B0(\key_mem[11][53] ), .B1(n4115), 
        .Y(n3220) );
  AO22X1 U2692 ( .A0(n4151), .A1(n667), .B0(\key_mem[9][53] ), .B1(n4160), .Y(
        n2964) );
  AO22X1 U2693 ( .A0(n4207), .A1(n667), .B0(\key_mem[7][53] ), .B1(n4215), .Y(
        n2708) );
  AO22X1 U2694 ( .A0(n4263), .A1(n667), .B0(\key_mem[5][53] ), .B1(n4280), .Y(
        n2452) );
  AO22X1 U2695 ( .A0(n4319), .A1(n667), .B0(\key_mem[3][53] ), .B1(n4341), .Y(
        n2196) );
  AO22X1 U2696 ( .A0(n4039), .A1(n1480), .B0(\key_mem[13][55] ), .B1(n4056), 
        .Y(n3474) );
  AO22X1 U2697 ( .A0(n4095), .A1(n665), .B0(\key_mem[11][55] ), .B1(n4107), 
        .Y(n3218) );
  AO22X1 U2698 ( .A0(n4151), .A1(n665), .B0(\key_mem[9][55] ), .B1(n4168), .Y(
        n2962) );
  AO22X1 U2699 ( .A0(n4207), .A1(n665), .B0(\key_mem[7][55] ), .B1(n4220), .Y(
        n2706) );
  AO22X1 U2700 ( .A0(n4263), .A1(n665), .B0(\key_mem[5][55] ), .B1(n4280), .Y(
        n2450) );
  AO22X1 U2701 ( .A0(n4319), .A1(n665), .B0(\key_mem[3][55] ), .B1(n4339), .Y(
        n2194) );
  AO22X1 U2702 ( .A0(n4040), .A1(n1490), .B0(\key_mem[13][65] ), .B1(n739), 
        .Y(n3464) );
  AO22X1 U2703 ( .A0(n4096), .A1(n655), .B0(\key_mem[11][65] ), .B1(n4113), 
        .Y(n3208) );
  AO22X1 U2704 ( .A0(n4152), .A1(n655), .B0(\key_mem[9][65] ), .B1(n4166), .Y(
        n2952) );
  AO22X1 U2705 ( .A0(n4208), .A1(n655), .B0(\key_mem[7][65] ), .B1(n4228), .Y(
        n2696) );
  AO22X1 U2706 ( .A0(n4264), .A1(n655), .B0(\key_mem[5][65] ), .B1(n4279), .Y(
        n2440) );
  AO22X1 U2707 ( .A0(n4320), .A1(n655), .B0(\key_mem[3][65] ), .B1(n4334), .Y(
        n2184) );
  AO22X1 U2708 ( .A0(n4040), .A1(n1491), .B0(\key_mem[13][66] ), .B1(n4059), 
        .Y(n3463) );
  AO22X1 U2709 ( .A0(n4096), .A1(n654), .B0(\key_mem[11][66] ), .B1(n4111), 
        .Y(n3207) );
  AO22X1 U2710 ( .A0(n4152), .A1(n654), .B0(\key_mem[9][66] ), .B1(n4165), .Y(
        n2951) );
  AO22X1 U2711 ( .A0(n4208), .A1(n654), .B0(\key_mem[7][66] ), .B1(n4227), .Y(
        n2695) );
  AO22X1 U2712 ( .A0(n4264), .A1(n654), .B0(\key_mem[5][66] ), .B1(n4272), .Y(
        n2439) );
  AO22X1 U2713 ( .A0(n4320), .A1(n654), .B0(\key_mem[3][66] ), .B1(n4341), .Y(
        n2183) );
  AO22X1 U2714 ( .A0(n4040), .A1(n1492), .B0(\key_mem[13][67] ), .B1(n4060), 
        .Y(n3462) );
  AO22X1 U2715 ( .A0(n4096), .A1(n653), .B0(\key_mem[11][67] ), .B1(n4112), 
        .Y(n3206) );
  AO22X1 U2716 ( .A0(n4152), .A1(n653), .B0(\key_mem[9][67] ), .B1(n4159), .Y(
        n2950) );
  AO22X1 U2717 ( .A0(n4208), .A1(n653), .B0(\key_mem[7][67] ), .B1(n4229), .Y(
        n2694) );
  AO22X1 U2718 ( .A0(n4264), .A1(n653), .B0(\key_mem[5][67] ), .B1(n4278), .Y(
        n2438) );
  AO22X1 U2719 ( .A0(n4320), .A1(n653), .B0(\key_mem[3][67] ), .B1(n4337), .Y(
        n2182) );
  AO22X1 U2720 ( .A0(n4040), .A1(n1493), .B0(\key_mem[13][68] ), .B1(n4061), 
        .Y(n3461) );
  AO22X1 U2721 ( .A0(n4096), .A1(n652), .B0(\key_mem[11][68] ), .B1(n737), .Y(
        n3205) );
  AO22X1 U2722 ( .A0(n4152), .A1(n652), .B0(\key_mem[9][68] ), .B1(n4160), .Y(
        n2949) );
  AO22X1 U2723 ( .A0(n4208), .A1(n652), .B0(\key_mem[7][68] ), .B1(n4229), .Y(
        n2693) );
  AO22X1 U2724 ( .A0(n4264), .A1(n652), .B0(\key_mem[5][68] ), .B1(n4271), .Y(
        n2437) );
  AO22X1 U2725 ( .A0(n4320), .A1(n652), .B0(\key_mem[3][68] ), .B1(n4328), .Y(
        n2181) );
  AO22X1 U2726 ( .A0(n4040), .A1(n1494), .B0(\key_mem[13][69] ), .B1(n4049), 
        .Y(n3460) );
  AO22X1 U2727 ( .A0(n4096), .A1(n651), .B0(\key_mem[11][69] ), .B1(n737), .Y(
        n3204) );
  AO22X1 U2728 ( .A0(n4152), .A1(n651), .B0(\key_mem[9][69] ), .B1(n4161), .Y(
        n2948) );
  AO22X1 U2729 ( .A0(n4208), .A1(n651), .B0(\key_mem[7][69] ), .B1(n4229), .Y(
        n2692) );
  AO22X1 U2730 ( .A0(n4264), .A1(n651), .B0(\key_mem[5][69] ), .B1(n4276), .Y(
        n2436) );
  AO22X1 U2731 ( .A0(n4320), .A1(n651), .B0(\key_mem[3][69] ), .B1(n4334), .Y(
        n2180) );
  AO22X1 U2732 ( .A0(n4041), .A1(n1496), .B0(\key_mem[13][71] ), .B1(n4056), 
        .Y(n3458) );
  AO22X1 U2733 ( .A0(n4097), .A1(n649), .B0(\key_mem[11][71] ), .B1(n737), .Y(
        n3202) );
  AO22X1 U2734 ( .A0(n4153), .A1(n649), .B0(\key_mem[9][71] ), .B1(n4164), .Y(
        n2946) );
  AO22X1 U2735 ( .A0(n4209), .A1(n649), .B0(\key_mem[7][71] ), .B1(n4229), .Y(
        n2690) );
  AO22X1 U2736 ( .A0(n4265), .A1(n649), .B0(\key_mem[5][71] ), .B1(n4273), .Y(
        n2434) );
  AO22X1 U2737 ( .A0(n4321), .A1(n649), .B0(\key_mem[3][71] ), .B1(n4339), .Y(
        n2178) );
  AO22X1 U2738 ( .A0(n4041), .A1(n1499), .B0(\key_mem[13][74] ), .B1(n4058), 
        .Y(n3455) );
  AO22X1 U2739 ( .A0(n4097), .A1(n646), .B0(\key_mem[11][74] ), .B1(n4108), 
        .Y(n3199) );
  AO22X1 U2740 ( .A0(n4153), .A1(n646), .B0(\key_mem[9][74] ), .B1(n4161), .Y(
        n2943) );
  AO22X1 U2741 ( .A0(n4209), .A1(n646), .B0(\key_mem[7][74] ), .B1(n4226), .Y(
        n2687) );
  AO22X1 U2742 ( .A0(n4265), .A1(n646), .B0(\key_mem[5][74] ), .B1(n4273), .Y(
        n2431) );
  AO22X1 U2743 ( .A0(n4321), .A1(n646), .B0(\key_mem[3][74] ), .B1(n4327), .Y(
        n2175) );
  AO22X1 U2744 ( .A0(n4041), .A1(n1502), .B0(\key_mem[13][77] ), .B1(n4056), 
        .Y(n3452) );
  AO22X1 U2745 ( .A0(n4097), .A1(n643), .B0(\key_mem[11][77] ), .B1(n4106), 
        .Y(n3196) );
  AO22X1 U2746 ( .A0(n4153), .A1(n643), .B0(\key_mem[9][77] ), .B1(n4164), .Y(
        n2940) );
  AO22X1 U2747 ( .A0(n4209), .A1(n643), .B0(\key_mem[7][77] ), .B1(n4218), .Y(
        n2684) );
  AO22X1 U2748 ( .A0(n4265), .A1(n643), .B0(\key_mem[5][77] ), .B1(n4274), .Y(
        n2428) );
  AO22X1 U2749 ( .A0(n4321), .A1(n643), .B0(\key_mem[3][77] ), .B1(n4328), .Y(
        n2172) );
  AO22X1 U2750 ( .A0(n4041), .A1(n1504), .B0(\key_mem[13][79] ), .B1(n4048), 
        .Y(n3450) );
  AO22X1 U2751 ( .A0(n4097), .A1(n641), .B0(\key_mem[11][79] ), .B1(n4108), 
        .Y(n3194) );
  AO22X1 U2752 ( .A0(n4153), .A1(n641), .B0(\key_mem[9][79] ), .B1(n4162), .Y(
        n2938) );
  AO22X1 U2753 ( .A0(n4209), .A1(n641), .B0(\key_mem[7][79] ), .B1(n4217), .Y(
        n2682) );
  AO22X1 U2754 ( .A0(n4265), .A1(n641), .B0(\key_mem[5][79] ), .B1(n4276), .Y(
        n2426) );
  AO22X1 U2755 ( .A0(n4321), .A1(n641), .B0(\key_mem[3][79] ), .B1(n4335), .Y(
        n2170) );
  AO22X1 U2756 ( .A0(n4042), .A1(n1506), .B0(\key_mem[13][81] ), .B1(n4047), 
        .Y(n3448) );
  AO22X1 U2757 ( .A0(n4098), .A1(n639), .B0(\key_mem[11][81] ), .B1(n4113), 
        .Y(n3192) );
  AO22X1 U2758 ( .A0(n4154), .A1(n639), .B0(\key_mem[9][81] ), .B1(n4163), .Y(
        n2936) );
  AO22X1 U2759 ( .A0(n4210), .A1(n639), .B0(\key_mem[7][81] ), .B1(n4226), .Y(
        n2680) );
  AO22X1 U2760 ( .A0(n4266), .A1(n639), .B0(\key_mem[5][81] ), .B1(n4275), .Y(
        n2424) );
  AO22X1 U2761 ( .A0(n4322), .A1(n639), .B0(\key_mem[3][81] ), .B1(n4334), .Y(
        n2168) );
  AO22X1 U2762 ( .A0(n4042), .A1(n1507), .B0(\key_mem[13][82] ), .B1(n4049), 
        .Y(n3447) );
  AO22X1 U2763 ( .A0(n4098), .A1(n638), .B0(\key_mem[11][82] ), .B1(n4112), 
        .Y(n3191) );
  AO22X1 U2764 ( .A0(n4154), .A1(n638), .B0(\key_mem[9][82] ), .B1(n4167), .Y(
        n2935) );
  AO22X1 U2765 ( .A0(n4210), .A1(n638), .B0(\key_mem[7][82] ), .B1(n4229), .Y(
        n2679) );
  AO22X1 U2766 ( .A0(n4266), .A1(n638), .B0(\key_mem[5][82] ), .B1(n4277), .Y(
        n2423) );
  AO22X1 U2767 ( .A0(n4322), .A1(n638), .B0(\key_mem[3][82] ), .B1(n4333), .Y(
        n2167) );
  AO22X1 U2768 ( .A0(n4042), .A1(n1509), .B0(\key_mem[13][84] ), .B1(n4058), 
        .Y(n3445) );
  AO22X1 U2769 ( .A0(n4098), .A1(n636), .B0(\key_mem[11][84] ), .B1(n4113), 
        .Y(n3189) );
  AO22X1 U2770 ( .A0(n4154), .A1(n636), .B0(\key_mem[9][84] ), .B1(n4161), .Y(
        n2933) );
  AO22X1 U2771 ( .A0(n4210), .A1(n636), .B0(\key_mem[7][84] ), .B1(n4216), .Y(
        n2677) );
  AO22X1 U2772 ( .A0(n4266), .A1(n636), .B0(\key_mem[5][84] ), .B1(n4273), .Y(
        n2421) );
  AO22X1 U2773 ( .A0(n4322), .A1(n636), .B0(\key_mem[3][84] ), .B1(n725), .Y(
        n2165) );
  AO22X1 U2774 ( .A0(n4042), .A1(n1510), .B0(\key_mem[13][85] ), .B1(n4059), 
        .Y(n3444) );
  AO22X1 U2775 ( .A0(n4098), .A1(n635), .B0(\key_mem[11][85] ), .B1(n4114), 
        .Y(n3188) );
  AO22X1 U2776 ( .A0(n4154), .A1(n635), .B0(\key_mem[9][85] ), .B1(n4167), .Y(
        n2932) );
  AO22X1 U2777 ( .A0(n4210), .A1(n635), .B0(\key_mem[7][85] ), .B1(n4227), .Y(
        n2676) );
  AO22X1 U2778 ( .A0(n4266), .A1(n635), .B0(\key_mem[5][85] ), .B1(n4272), .Y(
        n2420) );
  AO22X1 U2779 ( .A0(n4322), .A1(n635), .B0(\key_mem[3][85] ), .B1(n725), .Y(
        n2164) );
  AO22X1 U2780 ( .A0(n4042), .A1(n1512), .B0(\key_mem[13][87] ), .B1(n4049), 
        .Y(n3442) );
  AO22X1 U2781 ( .A0(n4098), .A1(n633), .B0(\key_mem[11][87] ), .B1(n4104), 
        .Y(n3186) );
  AO22X1 U2782 ( .A0(n4154), .A1(n633), .B0(\key_mem[9][87] ), .B1(n4159), .Y(
        n2930) );
  AO22X1 U2783 ( .A0(n4210), .A1(n633), .B0(\key_mem[7][87] ), .B1(n4220), .Y(
        n2674) );
  AO22X1 U2784 ( .A0(n4266), .A1(n633), .B0(\key_mem[5][87] ), .B1(n4271), .Y(
        n2418) );
  AO22X1 U2785 ( .A0(n4322), .A1(n633), .B0(\key_mem[3][87] ), .B1(n4327), .Y(
        n2162) );
  AO22X1 U2786 ( .A0(n4043), .A1(n1522), .B0(\key_mem[13][97] ), .B1(n4057), 
        .Y(n3432) );
  AO22X1 U2787 ( .A0(n4099), .A1(n623), .B0(\key_mem[11][97] ), .B1(n4114), 
        .Y(n3176) );
  AO22X1 U2788 ( .A0(n4155), .A1(n623), .B0(\key_mem[9][97] ), .B1(n4169), .Y(
        n2920) );
  AO22X1 U2789 ( .A0(n4211), .A1(n623), .B0(\key_mem[7][97] ), .B1(n4216), .Y(
        n2664) );
  AO22X1 U2790 ( .A0(n4267), .A1(n623), .B0(\key_mem[5][97] ), .B1(n4281), .Y(
        n2408) );
  AO22X1 U2791 ( .A0(n4323), .A1(n623), .B0(\key_mem[3][97] ), .B1(n4338), .Y(
        n2152) );
  AO22X1 U2792 ( .A0(n4043), .A1(n1523), .B0(\key_mem[13][98] ), .B1(n4057), 
        .Y(n3431) );
  AO22X1 U2793 ( .A0(n4099), .A1(n622), .B0(\key_mem[11][98] ), .B1(n4108), 
        .Y(n3175) );
  AO22X1 U2794 ( .A0(n4155), .A1(n622), .B0(\key_mem[9][98] ), .B1(n4168), .Y(
        n2919) );
  AO22X1 U2795 ( .A0(n4211), .A1(n622), .B0(\key_mem[7][98] ), .B1(n4217), .Y(
        n2663) );
  AO22X1 U2796 ( .A0(n4267), .A1(n622), .B0(\key_mem[5][98] ), .B1(n4280), .Y(
        n2407) );
  AO22X1 U2797 ( .A0(n4323), .A1(n622), .B0(\key_mem[3][98] ), .B1(n4341), .Y(
        n2151) );
  AO22X1 U2798 ( .A0(n4043), .A1(n1524), .B0(\key_mem[13][99] ), .B1(n4057), 
        .Y(n3430) );
  AO22X1 U2799 ( .A0(n4099), .A1(n621), .B0(\key_mem[11][99] ), .B1(n4106), 
        .Y(n3174) );
  AO22X1 U2800 ( .A0(n4155), .A1(n621), .B0(\key_mem[9][99] ), .B1(n4170), .Y(
        n2918) );
  AO22X1 U2801 ( .A0(n4211), .A1(n621), .B0(\key_mem[7][99] ), .B1(n4226), .Y(
        n2662) );
  AO22X1 U2802 ( .A0(n4267), .A1(n621), .B0(\key_mem[5][99] ), .B1(n4282), .Y(
        n2406) );
  AO22X1 U2803 ( .A0(n4323), .A1(n621), .B0(\key_mem[3][99] ), .B1(n4339), .Y(
        n2150) );
  AO22X1 U2804 ( .A0(n4044), .A1(n1525), .B0(\key_mem[13][100] ), .B1(n4057), 
        .Y(n3429) );
  AO22X1 U2805 ( .A0(n4100), .A1(n620), .B0(\key_mem[11][100] ), .B1(n4104), 
        .Y(n3173) );
  AO22X1 U2806 ( .A0(n4156), .A1(n620), .B0(\key_mem[9][100] ), .B1(n4169), 
        .Y(n2917) );
  AO22X1 U2807 ( .A0(n4212), .A1(n620), .B0(\key_mem[7][100] ), .B1(n4216), 
        .Y(n2661) );
  AO22X1 U2808 ( .A0(n4268), .A1(n620), .B0(\key_mem[5][100] ), .B1(n4281), 
        .Y(n2405) );
  AO22X1 U2809 ( .A0(n4324), .A1(n620), .B0(\key_mem[3][100] ), .B1(n4340), 
        .Y(n2149) );
  AO22X1 U2810 ( .A0(n4044), .A1(n1526), .B0(\key_mem[13][101] ), .B1(n4057), 
        .Y(n3428) );
  AO22X1 U2811 ( .A0(n4100), .A1(n619), .B0(\key_mem[11][101] ), .B1(n4103), 
        .Y(n3172) );
  AO22X1 U2812 ( .A0(n4156), .A1(n619), .B0(\key_mem[9][101] ), .B1(n4168), 
        .Y(n2916) );
  AO22X1 U2813 ( .A0(n4212), .A1(n619), .B0(\key_mem[7][101] ), .B1(n4215), 
        .Y(n2660) );
  AO22X1 U2814 ( .A0(n4268), .A1(n619), .B0(\key_mem[5][101] ), .B1(n4280), 
        .Y(n2404) );
  AO22X1 U2815 ( .A0(n4324), .A1(n619), .B0(\key_mem[3][101] ), .B1(n4331), 
        .Y(n2148) );
  AO22X1 U2816 ( .A0(n4044), .A1(n1528), .B0(\key_mem[13][103] ), .B1(n4056), 
        .Y(n3426) );
  AO22X1 U2817 ( .A0(n4100), .A1(n617), .B0(\key_mem[11][103] ), .B1(n4110), 
        .Y(n3170) );
  AO22X1 U2818 ( .A0(n4156), .A1(n617), .B0(\key_mem[9][103] ), .B1(n4168), 
        .Y(n2914) );
  AO22X1 U2819 ( .A0(n4212), .A1(n617), .B0(\key_mem[7][103] ), .B1(n4224), 
        .Y(n2658) );
  AO22X1 U2820 ( .A0(n4268), .A1(n617), .B0(\key_mem[5][103] ), .B1(n4280), 
        .Y(n2402) );
  AO22X1 U2821 ( .A0(n4324), .A1(n617), .B0(\key_mem[3][103] ), .B1(n4336), 
        .Y(n2146) );
  AO22X1 U2822 ( .A0(n4044), .A1(n1530), .B0(\key_mem[13][105] ), .B1(n4055), 
        .Y(n3424) );
  AO22X1 U2823 ( .A0(n4100), .A1(n615), .B0(\key_mem[11][105] ), .B1(n4115), 
        .Y(n3168) );
  AO22X1 U2824 ( .A0(n4156), .A1(n615), .B0(\key_mem[9][105] ), .B1(n4161), 
        .Y(n2912) );
  AO22X1 U2825 ( .A0(n4212), .A1(n615), .B0(\key_mem[7][105] ), .B1(n4224), 
        .Y(n2656) );
  AO22X1 U2826 ( .A0(n4268), .A1(n615), .B0(\key_mem[5][105] ), .B1(n4273), 
        .Y(n2400) );
  AO22X1 U2827 ( .A0(n4324), .A1(n615), .B0(\key_mem[3][105] ), .B1(n4336), 
        .Y(n2144) );
  AO22X1 U2828 ( .A0(n4044), .A1(n1531), .B0(\key_mem[13][106] ), .B1(n4049), 
        .Y(n3423) );
  AO22X1 U2829 ( .A0(n4100), .A1(n614), .B0(\key_mem[11][106] ), .B1(n4103), 
        .Y(n3167) );
  AO22X1 U2830 ( .A0(n4156), .A1(n614), .B0(\key_mem[9][106] ), .B1(n4159), 
        .Y(n2911) );
  AO22X1 U2831 ( .A0(n4212), .A1(n614), .B0(\key_mem[7][106] ), .B1(n4224), 
        .Y(n2655) );
  AO22X1 U2832 ( .A0(n4268), .A1(n614), .B0(\key_mem[5][106] ), .B1(n4272), 
        .Y(n2399) );
  AO22X1 U2833 ( .A0(n4324), .A1(n614), .B0(\key_mem[3][106] ), .B1(n4336), 
        .Y(n2143) );
  AO22X1 U2834 ( .A0(n4044), .A1(n1533), .B0(\key_mem[13][108] ), .B1(n4054), 
        .Y(n3421) );
  AO22X1 U2835 ( .A0(n4100), .A1(n612), .B0(\key_mem[11][108] ), .B1(n4105), 
        .Y(n3165) );
  AO22X1 U2836 ( .A0(n4156), .A1(n612), .B0(\key_mem[9][108] ), .B1(n4160), 
        .Y(n2909) );
  AO22X1 U2837 ( .A0(n4212), .A1(n612), .B0(\key_mem[7][108] ), .B1(n4224), 
        .Y(n2653) );
  AO22X1 U2838 ( .A0(n4268), .A1(n612), .B0(\key_mem[5][108] ), .B1(n4271), 
        .Y(n2397) );
  AO22X1 U2839 ( .A0(n4324), .A1(n612), .B0(\key_mem[3][108] ), .B1(n4336), 
        .Y(n2141) );
  AO22X1 U2840 ( .A0(n4044), .A1(n1534), .B0(\key_mem[13][109] ), .B1(n4047), 
        .Y(n3420) );
  AO22X1 U2841 ( .A0(n4100), .A1(n611), .B0(\key_mem[11][109] ), .B1(n4114), 
        .Y(n3164) );
  AO22X1 U2842 ( .A0(n4156), .A1(n611), .B0(\key_mem[9][109] ), .B1(n4164), 
        .Y(n2908) );
  AO22X1 U2843 ( .A0(n4212), .A1(n611), .B0(\key_mem[7][109] ), .B1(n4224), 
        .Y(n2652) );
  AO22X1 U2844 ( .A0(n4268), .A1(n611), .B0(\key_mem[5][109] ), .B1(n4276), 
        .Y(n2396) );
  AO22X1 U2845 ( .A0(n4324), .A1(n611), .B0(\key_mem[3][109] ), .B1(n4336), 
        .Y(n2140) );
  AO22X1 U2846 ( .A0(n4045), .A1(n1536), .B0(\key_mem[13][111] ), .B1(n4048), 
        .Y(n3418) );
  AO22X1 U2847 ( .A0(n4101), .A1(n609), .B0(\key_mem[11][111] ), .B1(n4113), 
        .Y(n3162) );
  AO22X1 U2848 ( .A0(n4157), .A1(n609), .B0(\key_mem[9][111] ), .B1(n4163), 
        .Y(n2906) );
  AO22X1 U2849 ( .A0(n4213), .A1(n609), .B0(\key_mem[7][111] ), .B1(n4224), 
        .Y(n2650) );
  AO22X1 U2850 ( .A0(n4269), .A1(n609), .B0(\key_mem[5][111] ), .B1(n4275), 
        .Y(n2394) );
  AO22X1 U2851 ( .A0(n4325), .A1(n609), .B0(\key_mem[3][111] ), .B1(n4336), 
        .Y(n2138) );
  AO22X1 U2852 ( .A0(n4045), .A1(n1537), .B0(\key_mem[13][112] ), .B1(n4051), 
        .Y(n3417) );
  AO22X1 U2853 ( .A0(n4101), .A1(n608), .B0(\key_mem[11][112] ), .B1(n4112), 
        .Y(n3161) );
  AO22X1 U2854 ( .A0(n4157), .A1(n608), .B0(\key_mem[9][112] ), .B1(n4162), 
        .Y(n2905) );
  AO22X1 U2855 ( .A0(n4213), .A1(n608), .B0(\key_mem[7][112] ), .B1(n4224), 
        .Y(n2649) );
  AO22X1 U2856 ( .A0(n4269), .A1(n608), .B0(\key_mem[5][112] ), .B1(n4274), 
        .Y(n2393) );
  AO22X1 U2857 ( .A0(n4325), .A1(n608), .B0(\key_mem[3][112] ), .B1(n4336), 
        .Y(n2137) );
  AO22X1 U2858 ( .A0(n4045), .A1(n1538), .B0(\key_mem[13][113] ), .B1(n4050), 
        .Y(n3416) );
  AO22X1 U2859 ( .A0(n4101), .A1(n607), .B0(\key_mem[11][113] ), .B1(n4106), 
        .Y(n3160) );
  AO22X1 U2860 ( .A0(n4157), .A1(n607), .B0(\key_mem[9][113] ), .B1(n4164), 
        .Y(n2904) );
  AO22X1 U2861 ( .A0(n4213), .A1(n607), .B0(\key_mem[7][113] ), .B1(n4225), 
        .Y(n2648) );
  AO22X1 U2862 ( .A0(n4269), .A1(n607), .B0(\key_mem[5][113] ), .B1(n4276), 
        .Y(n2392) );
  AO22X1 U2863 ( .A0(n4325), .A1(n607), .B0(\key_mem[3][113] ), .B1(n4329), 
        .Y(n2136) );
  AO22X1 U2864 ( .A0(n4045), .A1(n1539), .B0(\key_mem[13][114] ), .B1(n4049), 
        .Y(n3415) );
  AO22X1 U2865 ( .A0(n4101), .A1(n606), .B0(\key_mem[11][114] ), .B1(n4107), 
        .Y(n3159) );
  AO22X1 U2866 ( .A0(n4157), .A1(n606), .B0(\key_mem[9][114] ), .B1(n4163), 
        .Y(n2903) );
  AO22X1 U2867 ( .A0(n4213), .A1(n606), .B0(\key_mem[7][114] ), .B1(n4225), 
        .Y(n2647) );
  AO22X1 U2868 ( .A0(n4269), .A1(n606), .B0(\key_mem[5][114] ), .B1(n4275), 
        .Y(n2391) );
  AO22X1 U2869 ( .A0(n4325), .A1(n606), .B0(\key_mem[3][114] ), .B1(n4327), 
        .Y(n2135) );
  AO22X1 U2870 ( .A0(n4045), .A1(n1541), .B0(\key_mem[13][116] ), .B1(n4053), 
        .Y(n3413) );
  AO22X1 U2871 ( .A0(n4101), .A1(n604), .B0(\key_mem[11][116] ), .B1(n4114), 
        .Y(n3157) );
  AO22X1 U2872 ( .A0(n4157), .A1(n604), .B0(\key_mem[9][116] ), .B1(n4162), 
        .Y(n2901) );
  AO22X1 U2873 ( .A0(n4213), .A1(n604), .B0(\key_mem[7][116] ), .B1(n4225), 
        .Y(n2645) );
  AO22X1 U2874 ( .A0(n4269), .A1(n604), .B0(\key_mem[5][116] ), .B1(n4274), 
        .Y(n2389) );
  AO22X1 U2875 ( .A0(n4325), .A1(n604), .B0(\key_mem[3][116] ), .B1(n4328), 
        .Y(n2133) );
  AO22X1 U2876 ( .A0(n4045), .A1(n1542), .B0(\key_mem[13][117] ), .B1(n4052), 
        .Y(n3412) );
  AO22X1 U2877 ( .A0(n4101), .A1(n603), .B0(\key_mem[11][117] ), .B1(n4113), 
        .Y(n3156) );
  AO22X1 U2878 ( .A0(n4157), .A1(n603), .B0(\key_mem[9][117] ), .B1(n4167), 
        .Y(n2900) );
  AO22X1 U2879 ( .A0(n4213), .A1(n603), .B0(\key_mem[7][117] ), .B1(n4225), 
        .Y(n2644) );
  AO22X1 U2880 ( .A0(n4269), .A1(n603), .B0(\key_mem[5][117] ), .B1(n4279), 
        .Y(n2388) );
  AO22X1 U2881 ( .A0(n4325), .A1(n603), .B0(\key_mem[3][117] ), .B1(n4334), 
        .Y(n2132) );
  AO22X1 U2882 ( .A0(n4045), .A1(n1543), .B0(\key_mem[13][118] ), .B1(n4051), 
        .Y(n3411) );
  AO22X1 U2883 ( .A0(n4101), .A1(n602), .B0(\key_mem[11][118] ), .B1(n4112), 
        .Y(n3155) );
  AO22X1 U2884 ( .A0(n4157), .A1(n602), .B0(\key_mem[9][118] ), .B1(n4166), 
        .Y(n2899) );
  AO22X1 U2885 ( .A0(n4213), .A1(n602), .B0(\key_mem[7][118] ), .B1(n4225), 
        .Y(n2643) );
  AO22X1 U2886 ( .A0(n4269), .A1(n602), .B0(\key_mem[5][118] ), .B1(n4278), 
        .Y(n2387) );
  AO22X1 U2887 ( .A0(n4325), .A1(n602), .B0(\key_mem[3][118] ), .B1(n4332), 
        .Y(n2131) );
  AO22X1 U2888 ( .A0(n4045), .A1(n1544), .B0(\key_mem[13][119] ), .B1(n4050), 
        .Y(n3410) );
  AO22X1 U2889 ( .A0(n4101), .A1(n601), .B0(\key_mem[11][119] ), .B1(n4104), 
        .Y(n3154) );
  AO22X1 U2890 ( .A0(n4157), .A1(n601), .B0(\key_mem[9][119] ), .B1(n4165), 
        .Y(n2898) );
  AO22X1 U2891 ( .A0(n4213), .A1(n601), .B0(\key_mem[7][119] ), .B1(n4225), 
        .Y(n2642) );
  AO22X1 U2892 ( .A0(n4269), .A1(n601), .B0(\key_mem[5][119] ), .B1(n4277), 
        .Y(n2386) );
  AO22X1 U2893 ( .A0(n4325), .A1(n601), .B0(\key_mem[3][119] ), .B1(n4333), 
        .Y(n2130) );
  AO22X1 U2894 ( .A0(n4008), .A1(n1450), .B0(\key_mem[14][25] ), .B1(n4030), 
        .Y(n3632) );
  AO22X1 U2895 ( .A0(n4064), .A1(n1450), .B0(\key_mem[12][25] ), .B1(n4086), 
        .Y(n3376) );
  AO22X1 U2896 ( .A0(n4120), .A1(n1450), .B0(\key_mem[10][25] ), .B1(n4144), 
        .Y(n3120) );
  AO22X1 U2897 ( .A0(n4176), .A1(n1450), .B0(\key_mem[8][25] ), .B1(n4200), 
        .Y(n2864) );
  AO22X1 U2898 ( .A0(n4233), .A1(n1450), .B0(\key_mem[6][25] ), .B1(n4251), 
        .Y(n2608) );
  AO22X1 U2899 ( .A0(n4288), .A1(n1450), .B0(\key_mem[4][25] ), .B1(n4309), 
        .Y(n2352) );
  AO22X1 U2900 ( .A0(n4344), .A1(n1450), .B0(\key_mem[2][25] ), .B1(n4361), 
        .Y(n2096) );
  AO22X1 U2901 ( .A0(n3957), .A1(n1450), .B0(\key_mem[0][25] ), .B1(n1728), 
        .Y(n1840) );
  AO22X1 U2902 ( .A0(n4011), .A1(n1482), .B0(\key_mem[14][57] ), .B1(n4028), 
        .Y(n3600) );
  AO22X1 U2903 ( .A0(n4067), .A1(n1482), .B0(\key_mem[12][57] ), .B1(n4082), 
        .Y(n3344) );
  AO22X1 U2904 ( .A0(n4123), .A1(n1482), .B0(\key_mem[10][57] ), .B1(n4145), 
        .Y(n3088) );
  AO22X1 U2905 ( .A0(n4179), .A1(n1482), .B0(\key_mem[8][57] ), .B1(n4201), 
        .Y(n2832) );
  AO22X1 U2906 ( .A0(n4236), .A1(n1482), .B0(\key_mem[6][57] ), .B1(n4230), 
        .Y(n2576) );
  AO22X1 U2907 ( .A0(n4291), .A1(n1482), .B0(\key_mem[4][57] ), .B1(n4311), 
        .Y(n2320) );
  AO22X1 U2908 ( .A0(n4347), .A1(n1482), .B0(\key_mem[2][57] ), .B1(n4360), 
        .Y(n2064) );
  AO22X1 U2909 ( .A0(n3954), .A1(n1482), .B0(\key_mem[0][57] ), .B1(n3929), 
        .Y(n1808) );
  AO22X1 U2910 ( .A0(n4014), .A1(n1514), .B0(\key_mem[14][89] ), .B1(n4028), 
        .Y(n3568) );
  AO22X1 U2911 ( .A0(n4070), .A1(n1514), .B0(\key_mem[12][89] ), .B1(n4081), 
        .Y(n3312) );
  AO22X1 U2912 ( .A0(n4126), .A1(n1514), .B0(\key_mem[10][89] ), .B1(n4140), 
        .Y(n3056) );
  AO22X1 U2913 ( .A0(n4182), .A1(n1514), .B0(\key_mem[8][89] ), .B1(n4196), 
        .Y(n2800) );
  AO22X1 U2914 ( .A0(n4239), .A1(n1514), .B0(\key_mem[6][89] ), .B1(n4245), 
        .Y(n2544) );
  AO22X1 U2915 ( .A0(n4294), .A1(n1514), .B0(\key_mem[4][89] ), .B1(n4306), 
        .Y(n2288) );
  AO22X1 U2916 ( .A0(n4350), .A1(n1514), .B0(\key_mem[2][89] ), .B1(n4357), 
        .Y(n2032) );
  AO22X1 U2917 ( .A0(n3951), .A1(n1514), .B0(\key_mem[0][89] ), .B1(n3932), 
        .Y(n1776) );
  AO22X1 U2918 ( .A0(n4018), .A1(n1546), .B0(\key_mem[14][121] ), .B1(n4033), 
        .Y(n3536) );
  AO22X1 U2919 ( .A0(n4074), .A1(n1546), .B0(\key_mem[12][121] ), .B1(n4085), 
        .Y(n3280) );
  AO22X1 U2920 ( .A0(n4130), .A1(n1546), .B0(\key_mem[10][121] ), .B1(n4140), 
        .Y(n3024) );
  AO22X1 U2921 ( .A0(n4186), .A1(n1546), .B0(\key_mem[8][121] ), .B1(n4196), 
        .Y(n2768) );
  AO22X1 U2922 ( .A0(n4243), .A1(n1546), .B0(\key_mem[6][121] ), .B1(n4254), 
        .Y(n2512) );
  AO22X1 U2923 ( .A0(n4298), .A1(n1546), .B0(\key_mem[4][121] ), .B1(n4308), 
        .Y(n2256) );
  AO22X1 U2924 ( .A0(n4354), .A1(n1546), .B0(\key_mem[2][121] ), .B1(n4365), 
        .Y(n2000) );
  AO22X1 U2925 ( .A0(n3962), .A1(n1546), .B0(\key_mem[0][121] ), .B1(n3934), 
        .Y(n1744) );
  AO22X1 U2926 ( .A0(n4008), .A1(n1453), .B0(\key_mem[14][28] ), .B1(n4031), 
        .Y(n3629) );
  AO22X1 U2927 ( .A0(n4064), .A1(n1453), .B0(\key_mem[12][28] ), .B1(n4089), 
        .Y(n3373) );
  AO22X1 U2928 ( .A0(n4120), .A1(n1453), .B0(\key_mem[10][28] ), .B1(n4139), 
        .Y(n3117) );
  AO22X1 U2929 ( .A0(n4176), .A1(n1453), .B0(\key_mem[8][28] ), .B1(n4195), 
        .Y(n2861) );
  AO22X1 U2930 ( .A0(n4233), .A1(n1453), .B0(\key_mem[6][28] ), .B1(n730), .Y(
        n2605) );
  AO22X1 U2931 ( .A0(n4288), .A1(n1453), .B0(\key_mem[4][28] ), .B1(n4303), 
        .Y(n2349) );
  AO22X1 U2932 ( .A0(n4344), .A1(n1453), .B0(\key_mem[2][28] ), .B1(n4365), 
        .Y(n2093) );
  AO22X1 U2933 ( .A0(n3957), .A1(n1453), .B0(\key_mem[0][28] ), .B1(n1728), 
        .Y(n1837) );
  AO22X1 U2934 ( .A0(n4012), .A1(n1485), .B0(\key_mem[14][60] ), .B1(n4027), 
        .Y(n3597) );
  AO22X1 U2935 ( .A0(n4068), .A1(n1485), .B0(\key_mem[12][60] ), .B1(n4081), 
        .Y(n3341) );
  AO22X1 U2936 ( .A0(n4124), .A1(n1485), .B0(\key_mem[10][60] ), .B1(n4135), 
        .Y(n3085) );
  AO22X1 U2937 ( .A0(n4180), .A1(n1485), .B0(\key_mem[8][60] ), .B1(n4191), 
        .Y(n2829) );
  AO22X1 U2938 ( .A0(n4237), .A1(n1485), .B0(\key_mem[6][60] ), .B1(n4248), 
        .Y(n2573) );
  AO22X1 U2939 ( .A0(n4292), .A1(n1485), .B0(\key_mem[4][60] ), .B1(n4312), 
        .Y(n2317) );
  AO22X1 U2940 ( .A0(n4348), .A1(n1485), .B0(\key_mem[2][60] ), .B1(n4356), 
        .Y(n2061) );
  AO22X1 U2941 ( .A0(n3954), .A1(n1485), .B0(\key_mem[0][60] ), .B1(n3929), 
        .Y(n1805) );
  AO22X1 U2942 ( .A0(n4015), .A1(n1517), .B0(\key_mem[14][92] ), .B1(n4027), 
        .Y(n3565) );
  AO22X1 U2943 ( .A0(n4071), .A1(n1517), .B0(\key_mem[12][92] ), .B1(n4080), 
        .Y(n3309) );
  AO22X1 U2944 ( .A0(n4127), .A1(n1517), .B0(\key_mem[10][92] ), .B1(n4141), 
        .Y(n3053) );
  AO22X1 U2945 ( .A0(n4183), .A1(n1517), .B0(\key_mem[8][92] ), .B1(n4197), 
        .Y(n2797) );
  AO22X1 U2946 ( .A0(n4240), .A1(n1517), .B0(\key_mem[6][92] ), .B1(n4245), 
        .Y(n2541) );
  AO22X1 U2947 ( .A0(n4295), .A1(n1517), .B0(\key_mem[4][92] ), .B1(n4307), 
        .Y(n2285) );
  AO22X1 U2948 ( .A0(n4351), .A1(n1517), .B0(\key_mem[2][92] ), .B1(n4356), 
        .Y(n2029) );
  AO22X1 U2949 ( .A0(n3951), .A1(n1517), .B0(\key_mem[0][92] ), .B1(n3932), 
        .Y(n1773) );
  AO22X1 U2950 ( .A0(n4018), .A1(n1549), .B0(\key_mem[14][124] ), .B1(n4027), 
        .Y(n3533) );
  AO22X1 U2951 ( .A0(n4074), .A1(n1549), .B0(\key_mem[12][124] ), .B1(n4086), 
        .Y(n3277) );
  AO22X1 U2952 ( .A0(n4130), .A1(n1549), .B0(\key_mem[10][124] ), .B1(n4135), 
        .Y(n3021) );
  AO22X1 U2953 ( .A0(n4186), .A1(n1549), .B0(\key_mem[8][124] ), .B1(n4191), 
        .Y(n2765) );
  AO22X1 U2954 ( .A0(n4243), .A1(n1549), .B0(\key_mem[6][124] ), .B1(n4256), 
        .Y(n2509) );
  AO22X1 U2955 ( .A0(n4298), .A1(n1549), .B0(\key_mem[4][124] ), .B1(n4304), 
        .Y(n2253) );
  AO22X1 U2956 ( .A0(n4354), .A1(n1549), .B0(\key_mem[2][124] ), .B1(n4356), 
        .Y(n1997) );
  AO22X1 U2957 ( .A0(n3960), .A1(n1549), .B0(\key_mem[0][124] ), .B1(n3934), 
        .Y(n1741) );
  AO22X1 U2958 ( .A0(n4008), .A1(n1454), .B0(\key_mem[14][29] ), .B1(n4032), 
        .Y(n3628) );
  AO22X1 U2959 ( .A0(n4064), .A1(n1454), .B0(\key_mem[12][29] ), .B1(n4088), 
        .Y(n3372) );
  AO22X1 U2960 ( .A0(n4120), .A1(n1454), .B0(\key_mem[10][29] ), .B1(n4143), 
        .Y(n3116) );
  AO22X1 U2961 ( .A0(n4176), .A1(n1454), .B0(\key_mem[8][29] ), .B1(n4199), 
        .Y(n2860) );
  AO22X1 U2962 ( .A0(n4233), .A1(n1454), .B0(\key_mem[6][29] ), .B1(n4255), 
        .Y(n2604) );
  AO22X1 U2963 ( .A0(n4288), .A1(n1454), .B0(\key_mem[4][29] ), .B1(n4308), 
        .Y(n2348) );
  AO22X1 U2964 ( .A0(n4344), .A1(n1454), .B0(\key_mem[2][29] ), .B1(n4364), 
        .Y(n2092) );
  AO22X1 U2965 ( .A0(n3957), .A1(n1454), .B0(\key_mem[0][29] ), .B1(n1728), 
        .Y(n1836) );
  AO22X1 U2966 ( .A0(n4012), .A1(n1486), .B0(\key_mem[14][61] ), .B1(n4029), 
        .Y(n3596) );
  AO22X1 U2967 ( .A0(n4068), .A1(n1486), .B0(\key_mem[12][61] ), .B1(n4077), 
        .Y(n3340) );
  AO22X1 U2968 ( .A0(n4124), .A1(n1486), .B0(\key_mem[10][61] ), .B1(n4142), 
        .Y(n3084) );
  AO22X1 U2969 ( .A0(n4180), .A1(n1486), .B0(\key_mem[8][61] ), .B1(n4198), 
        .Y(n2828) );
  AO22X1 U2970 ( .A0(n4237), .A1(n1486), .B0(\key_mem[6][61] ), .B1(n4249), 
        .Y(n2572) );
  AO22X1 U2971 ( .A0(n4292), .A1(n1486), .B0(\key_mem[4][61] ), .B1(n4304), 
        .Y(n2316) );
  AO22X1 U2972 ( .A0(n4348), .A1(n1486), .B0(\key_mem[2][61] ), .B1(n722), .Y(
        n2060) );
  AO22X1 U2973 ( .A0(n3954), .A1(n1486), .B0(\key_mem[0][61] ), .B1(n3930), 
        .Y(n1804) );
  AO22X1 U2974 ( .A0(n4015), .A1(n1518), .B0(\key_mem[14][93] ), .B1(n4025), 
        .Y(n3564) );
  AO22X1 U2975 ( .A0(n4071), .A1(n1518), .B0(\key_mem[12][93] ), .B1(n4086), 
        .Y(n3308) );
  AO22X1 U2976 ( .A0(n4127), .A1(n1518), .B0(\key_mem[10][93] ), .B1(n4140), 
        .Y(n3052) );
  AO22X1 U2977 ( .A0(n4183), .A1(n1518), .B0(\key_mem[8][93] ), .B1(n4196), 
        .Y(n2796) );
  AO22X1 U2978 ( .A0(n4240), .A1(n1518), .B0(\key_mem[6][93] ), .B1(n4245), 
        .Y(n2540) );
  AO22X1 U2979 ( .A0(n4295), .A1(n1518), .B0(\key_mem[4][93] ), .B1(n4307), 
        .Y(n2284) );
  AO22X1 U2980 ( .A0(n4351), .A1(n1518), .B0(\key_mem[2][93] ), .B1(n4365), 
        .Y(n2028) );
  AO22X1 U2981 ( .A0(n3950), .A1(n1518), .B0(\key_mem[0][93] ), .B1(n3932), 
        .Y(n1772) );
  AO22X1 U2982 ( .A0(n4018), .A1(n1550), .B0(\key_mem[14][125] ), .B1(n4029), 
        .Y(n3532) );
  AO22X1 U2983 ( .A0(n4074), .A1(n1550), .B0(\key_mem[12][125] ), .B1(n4088), 
        .Y(n3276) );
  AO22X1 U2984 ( .A0(n4130), .A1(n1550), .B0(\key_mem[10][125] ), .B1(n4134), 
        .Y(n3020) );
  AO22X1 U2985 ( .A0(n4186), .A1(n1550), .B0(\key_mem[8][125] ), .B1(n4190), 
        .Y(n2764) );
  AO22X1 U2986 ( .A0(n4243), .A1(n1550), .B0(\key_mem[6][125] ), .B1(n4230), 
        .Y(n2508) );
  AO22X1 U2987 ( .A0(n4298), .A1(n1550), .B0(\key_mem[4][125] ), .B1(n4303), 
        .Y(n2252) );
  AO22X1 U2988 ( .A0(n4354), .A1(n1550), .B0(\key_mem[2][125] ), .B1(n4355), 
        .Y(n1996) );
  AO22X1 U2989 ( .A0(n3963), .A1(n1550), .B0(\key_mem[0][125] ), .B1(n3934), 
        .Y(n1740) );
  AO22X1 U2990 ( .A0(n4009), .A1(n1455), .B0(\key_mem[14][30] ), .B1(n4033), 
        .Y(n3627) );
  AO22X1 U2991 ( .A0(n4065), .A1(n1455), .B0(\key_mem[12][30] ), .B1(n4083), 
        .Y(n3371) );
  AO22X1 U2992 ( .A0(n4121), .A1(n1455), .B0(\key_mem[10][30] ), .B1(n4144), 
        .Y(n3115) );
  AO22X1 U2993 ( .A0(n4177), .A1(n1455), .B0(\key_mem[8][30] ), .B1(n4200), 
        .Y(n2859) );
  AO22X1 U2994 ( .A0(n4234), .A1(n1455), .B0(\key_mem[6][30] ), .B1(n4255), 
        .Y(n2603) );
  AO22X1 U2995 ( .A0(n4289), .A1(n1455), .B0(\key_mem[4][30] ), .B1(n4310), 
        .Y(n2347) );
  AO22X1 U2996 ( .A0(n4345), .A1(n1455), .B0(\key_mem[2][30] ), .B1(n4363), 
        .Y(n2091) );
  AO22X1 U2997 ( .A0(n3957), .A1(n1455), .B0(\key_mem[0][30] ), .B1(n1728), 
        .Y(n1835) );
  AO22X1 U2998 ( .A0(n4012), .A1(n1487), .B0(\key_mem[14][62] ), .B1(n4030), 
        .Y(n3595) );
  AO22X1 U2999 ( .A0(n4068), .A1(n1487), .B0(\key_mem[12][62] ), .B1(n4080), 
        .Y(n3339) );
  AO22X1 U3000 ( .A0(n4124), .A1(n1487), .B0(\key_mem[10][62] ), .B1(n4141), 
        .Y(n3083) );
  AO22X1 U3001 ( .A0(n4180), .A1(n1487), .B0(\key_mem[8][62] ), .B1(n4197), 
        .Y(n2827) );
  AO22X1 U3002 ( .A0(n4237), .A1(n1487), .B0(\key_mem[6][62] ), .B1(n4251), 
        .Y(n2571) );
  AO22X1 U3003 ( .A0(n4292), .A1(n1487), .B0(\key_mem[4][62] ), .B1(n727), .Y(
        n2315) );
  AO22X1 U3004 ( .A0(n4348), .A1(n1487), .B0(\key_mem[2][62] ), .B1(n4367), 
        .Y(n2059) );
  AO22X1 U3005 ( .A0(n3954), .A1(n1487), .B0(\key_mem[0][62] ), .B1(n3930), 
        .Y(n1803) );
  AO22X1 U3006 ( .A0(n4015), .A1(n1519), .B0(\key_mem[14][94] ), .B1(n4023), 
        .Y(n3563) );
  AO22X1 U3007 ( .A0(n4071), .A1(n1519), .B0(\key_mem[12][94] ), .B1(n4080), 
        .Y(n3307) );
  AO22X1 U3008 ( .A0(n4127), .A1(n1519), .B0(\key_mem[10][94] ), .B1(n4142), 
        .Y(n3051) );
  AO22X1 U3009 ( .A0(n4183), .A1(n1519), .B0(\key_mem[8][94] ), .B1(n4198), 
        .Y(n2795) );
  AO22X1 U3010 ( .A0(n4240), .A1(n1519), .B0(\key_mem[6][94] ), .B1(n4253), 
        .Y(n2539) );
  AO22X1 U3011 ( .A0(n4295), .A1(n1519), .B0(\key_mem[4][94] ), .B1(n4305), 
        .Y(n2283) );
  AO22X1 U3012 ( .A0(n4351), .A1(n1519), .B0(\key_mem[2][94] ), .B1(n4365), 
        .Y(n2027) );
  AO22X1 U3013 ( .A0(n3950), .A1(n1519), .B0(\key_mem[0][94] ), .B1(n3932), 
        .Y(n1771) );
  AO22X1 U3014 ( .A0(n4018), .A1(n1551), .B0(\key_mem[14][126] ), .B1(n4019), 
        .Y(n3531) );
  AO22X1 U3015 ( .A0(n4074), .A1(n1551), .B0(\key_mem[12][126] ), .B1(n4089), 
        .Y(n3275) );
  AO22X1 U3016 ( .A0(n4130), .A1(n1551), .B0(\key_mem[10][126] ), .B1(n4133), 
        .Y(n3019) );
  AO22X1 U3017 ( .A0(n4186), .A1(n1551), .B0(\key_mem[8][126] ), .B1(n4189), 
        .Y(n2763) );
  AO22X1 U3018 ( .A0(n4243), .A1(n1551), .B0(\key_mem[6][126] ), .B1(n4230), 
        .Y(n2507) );
  AO22X1 U3019 ( .A0(n4298), .A1(n1551), .B0(\key_mem[4][126] ), .B1(n4302), 
        .Y(n2251) );
  AO22X1 U3020 ( .A0(n4354), .A1(n1551), .B0(\key_mem[2][126] ), .B1(n4360), 
        .Y(n1995) );
  AO22X1 U3021 ( .A0(n3963), .A1(n1551), .B0(\key_mem[0][126] ), .B1(n3934), 
        .Y(n1739) );
  AO22X1 U3022 ( .A0(n4008), .A1(n1452), .B0(\key_mem[14][27] ), .B1(n4021), 
        .Y(n3630) );
  AO22X1 U3023 ( .A0(n4064), .A1(n1452), .B0(\key_mem[12][27] ), .B1(n4089), 
        .Y(n3374) );
  AO22X1 U3024 ( .A0(n4120), .A1(n1452), .B0(\key_mem[10][27] ), .B1(n4145), 
        .Y(n3118) );
  AO22X1 U3025 ( .A0(n4176), .A1(n1452), .B0(\key_mem[8][27] ), .B1(n4201), 
        .Y(n2862) );
  AO22X1 U3026 ( .A0(n4233), .A1(n1452), .B0(\key_mem[6][27] ), .B1(n4256), 
        .Y(n2606) );
  AO22X1 U3027 ( .A0(n4288), .A1(n1452), .B0(\key_mem[4][27] ), .B1(n4299), 
        .Y(n2350) );
  AO22X1 U3028 ( .A0(n4344), .A1(n1452), .B0(\key_mem[2][27] ), .B1(n4362), 
        .Y(n2094) );
  AO22X1 U3029 ( .A0(n3957), .A1(n1452), .B0(\key_mem[0][27] ), .B1(n1728), 
        .Y(n1838) );
  AO22X1 U3030 ( .A0(n4011), .A1(n1484), .B0(\key_mem[14][59] ), .B1(n4028), 
        .Y(n3598) );
  AO22X1 U3031 ( .A0(n4067), .A1(n1484), .B0(\key_mem[12][59] ), .B1(n4079), 
        .Y(n3342) );
  AO22X1 U3032 ( .A0(n4123), .A1(n1484), .B0(\key_mem[10][59] ), .B1(n4136), 
        .Y(n3086) );
  AO22X1 U3033 ( .A0(n4179), .A1(n1484), .B0(\key_mem[8][59] ), .B1(n4192), 
        .Y(n2830) );
  AO22X1 U3034 ( .A0(n4236), .A1(n1484), .B0(\key_mem[6][59] ), .B1(n4246), 
        .Y(n2574) );
  AO22X1 U3035 ( .A0(n4291), .A1(n1484), .B0(\key_mem[4][59] ), .B1(n4311), 
        .Y(n2318) );
  AO22X1 U3036 ( .A0(n4347), .A1(n1484), .B0(\key_mem[2][59] ), .B1(n4368), 
        .Y(n2062) );
  AO22X1 U3037 ( .A0(n3954), .A1(n1484), .B0(\key_mem[0][59] ), .B1(n3929), 
        .Y(n1806) );
  AO22X1 U3038 ( .A0(n4015), .A1(n1516), .B0(\key_mem[14][91] ), .B1(n4029), 
        .Y(n3566) );
  AO22X1 U3039 ( .A0(n4071), .A1(n1516), .B0(\key_mem[12][91] ), .B1(n4078), 
        .Y(n3310) );
  AO22X1 U3040 ( .A0(n4127), .A1(n1516), .B0(\key_mem[10][91] ), .B1(n4140), 
        .Y(n3054) );
  AO22X1 U3041 ( .A0(n4183), .A1(n1516), .B0(\key_mem[8][91] ), .B1(n4196), 
        .Y(n2798) );
  AO22X1 U3042 ( .A0(n4240), .A1(n1516), .B0(\key_mem[6][91] ), .B1(n4253), 
        .Y(n2542) );
  AO22X1 U3043 ( .A0(n4295), .A1(n1516), .B0(\key_mem[4][91] ), .B1(n4305), 
        .Y(n2286) );
  AO22X1 U3044 ( .A0(n4351), .A1(n1516), .B0(\key_mem[2][91] ), .B1(n4355), 
        .Y(n2030) );
  AO22X1 U3045 ( .A0(n3951), .A1(n1516), .B0(\key_mem[0][91] ), .B1(n3932), 
        .Y(n1774) );
  AO22X1 U3046 ( .A0(n4018), .A1(n1548), .B0(\key_mem[14][123] ), .B1(n4026), 
        .Y(n3534) );
  AO22X1 U3047 ( .A0(n4074), .A1(n1548), .B0(\key_mem[12][123] ), .B1(n4075), 
        .Y(n3278) );
  AO22X1 U3048 ( .A0(n4130), .A1(n1548), .B0(\key_mem[10][123] ), .B1(n4131), 
        .Y(n3022) );
  AO22X1 U3049 ( .A0(n4186), .A1(n1548), .B0(\key_mem[8][123] ), .B1(n4187), 
        .Y(n2766) );
  AO22X1 U3050 ( .A0(n4243), .A1(n1548), .B0(\key_mem[6][123] ), .B1(n730), 
        .Y(n2510) );
  AO22X1 U3051 ( .A0(n4298), .A1(n1548), .B0(\key_mem[4][123] ), .B1(n4301), 
        .Y(n2254) );
  AO22X1 U3052 ( .A0(n4354), .A1(n1548), .B0(\key_mem[2][123] ), .B1(n4359), 
        .Y(n1998) );
  AO22X1 U3053 ( .A0(n3963), .A1(n1548), .B0(\key_mem[0][123] ), .B1(n3934), 
        .Y(n1742) );
  AO22X1 U3054 ( .A0(n4008), .A1(n1451), .B0(\key_mem[14][26] ), .B1(n4032), 
        .Y(n3631) );
  AO22X1 U3055 ( .A0(n4064), .A1(n1451), .B0(\key_mem[12][26] ), .B1(n4078), 
        .Y(n3375) );
  AO22X1 U3056 ( .A0(n4120), .A1(n1451), .B0(\key_mem[10][26] ), .B1(n4138), 
        .Y(n3119) );
  AO22X1 U3057 ( .A0(n4176), .A1(n1451), .B0(\key_mem[8][26] ), .B1(n4194), 
        .Y(n2863) );
  AO22X1 U3058 ( .A0(n4233), .A1(n1451), .B0(\key_mem[6][26] ), .B1(n4256), 
        .Y(n2607) );
  AO22X1 U3059 ( .A0(n4288), .A1(n1451), .B0(\key_mem[4][26] ), .B1(n4302), 
        .Y(n2351) );
  AO22X1 U3060 ( .A0(n4344), .A1(n1451), .B0(\key_mem[2][26] ), .B1(n4361), 
        .Y(n2095) );
  AO22X1 U3061 ( .A0(n3957), .A1(n1451), .B0(\key_mem[0][26] ), .B1(n1728), 
        .Y(n1839) );
  AO22X1 U3062 ( .A0(n4011), .A1(n1483), .B0(\key_mem[14][58] ), .B1(n4027), 
        .Y(n3599) );
  AO22X1 U3063 ( .A0(n4067), .A1(n1483), .B0(\key_mem[12][58] ), .B1(n4078), 
        .Y(n3343) );
  AO22X1 U3064 ( .A0(n4123), .A1(n1483), .B0(\key_mem[10][58] ), .B1(n4135), 
        .Y(n3087) );
  AO22X1 U3065 ( .A0(n4179), .A1(n1483), .B0(\key_mem[8][58] ), .B1(n4191), 
        .Y(n2831) );
  AO22X1 U3066 ( .A0(n4236), .A1(n1483), .B0(\key_mem[6][58] ), .B1(n4252), 
        .Y(n2575) );
  AO22X1 U3067 ( .A0(n4291), .A1(n1483), .B0(\key_mem[4][58] ), .B1(n4312), 
        .Y(n2319) );
  AO22X1 U3068 ( .A0(n4347), .A1(n1483), .B0(\key_mem[2][58] ), .B1(n4369), 
        .Y(n2063) );
  AO22X1 U3069 ( .A0(n3954), .A1(n1483), .B0(\key_mem[0][58] ), .B1(n3929), 
        .Y(n1807) );
  AO22X1 U3070 ( .A0(n4015), .A1(n1515), .B0(\key_mem[14][90] ), .B1(n4020), 
        .Y(n3567) );
  AO22X1 U3071 ( .A0(n4071), .A1(n1515), .B0(\key_mem[12][90] ), .B1(n4076), 
        .Y(n3311) );
  AO22X1 U3072 ( .A0(n4127), .A1(n1515), .B0(\key_mem[10][90] ), .B1(n4142), 
        .Y(n3055) );
  AO22X1 U3073 ( .A0(n4183), .A1(n1515), .B0(\key_mem[8][90] ), .B1(n4198), 
        .Y(n2799) );
  AO22X1 U3074 ( .A0(n4240), .A1(n1515), .B0(\key_mem[6][90] ), .B1(n4246), 
        .Y(n2543) );
  AO22X1 U3075 ( .A0(n4295), .A1(n1515), .B0(\key_mem[4][90] ), .B1(n4303), 
        .Y(n2287) );
  AO22X1 U3076 ( .A0(n4351), .A1(n1515), .B0(\key_mem[2][90] ), .B1(n4364), 
        .Y(n2031) );
  AO22X1 U3077 ( .A0(n3951), .A1(n1515), .B0(\key_mem[0][90] ), .B1(n3932), 
        .Y(n1775) );
  AO22X1 U3078 ( .A0(n4018), .A1(n1547), .B0(\key_mem[14][122] ), .B1(n4030), 
        .Y(n3535) );
  AO22X1 U3079 ( .A0(n4074), .A1(n1547), .B0(\key_mem[12][122] ), .B1(n4085), 
        .Y(n3279) );
  AO22X1 U3080 ( .A0(n4130), .A1(n1547), .B0(\key_mem[10][122] ), .B1(n4131), 
        .Y(n3023) );
  AO22X1 U3081 ( .A0(n4186), .A1(n1547), .B0(\key_mem[8][122] ), .B1(n4187), 
        .Y(n2767) );
  AO22X1 U3082 ( .A0(n4243), .A1(n1547), .B0(\key_mem[6][122] ), .B1(n4246), 
        .Y(n2511) );
  AO22X1 U3083 ( .A0(n4298), .A1(n1547), .B0(\key_mem[4][122] ), .B1(n4309), 
        .Y(n2255) );
  AO22X1 U3084 ( .A0(n4354), .A1(n1547), .B0(\key_mem[2][122] ), .B1(n4364), 
        .Y(n1999) );
  AO22X1 U3085 ( .A0(n3960), .A1(n1547), .B0(\key_mem[0][122] ), .B1(n3934), 
        .Y(n1743) );
  AO22X1 U3086 ( .A0(n4008), .A1(n1449), .B0(\key_mem[14][24] ), .B1(n4022), 
        .Y(n3633) );
  AO22X1 U3087 ( .A0(n4064), .A1(n1449), .B0(\key_mem[12][24] ), .B1(n4082), 
        .Y(n3377) );
  AO22X1 U3088 ( .A0(n4120), .A1(n1449), .B0(\key_mem[10][24] ), .B1(n4137), 
        .Y(n3121) );
  AO22X1 U3089 ( .A0(n4176), .A1(n1449), .B0(\key_mem[8][24] ), .B1(n4193), 
        .Y(n2865) );
  AO22X1 U3090 ( .A0(n4233), .A1(n1449), .B0(\key_mem[6][24] ), .B1(n4244), 
        .Y(n2609) );
  AO22X1 U3091 ( .A0(n4288), .A1(n1449), .B0(\key_mem[4][24] ), .B1(n4299), 
        .Y(n2353) );
  AO22X1 U3092 ( .A0(n4344), .A1(n1449), .B0(\key_mem[2][24] ), .B1(n4360), 
        .Y(n2097) );
  AO22X1 U3093 ( .A0(n3957), .A1(n1449), .B0(\key_mem[0][24] ), .B1(n1728), 
        .Y(n1841) );
  AO22X1 U3094 ( .A0(n4011), .A1(n1481), .B0(\key_mem[14][56] ), .B1(n4029), 
        .Y(n3601) );
  AO22X1 U3095 ( .A0(n4067), .A1(n1481), .B0(\key_mem[12][56] ), .B1(n4077), 
        .Y(n3345) );
  AO22X1 U3096 ( .A0(n4123), .A1(n1481), .B0(\key_mem[10][56] ), .B1(n4140), 
        .Y(n3089) );
  AO22X1 U3097 ( .A0(n4179), .A1(n1481), .B0(\key_mem[8][56] ), .B1(n4196), 
        .Y(n2833) );
  AO22X1 U3098 ( .A0(n4236), .A1(n1481), .B0(\key_mem[6][56] ), .B1(n4251), 
        .Y(n2577) );
  AO22X1 U3099 ( .A0(n4291), .A1(n1481), .B0(\key_mem[4][56] ), .B1(n4313), 
        .Y(n2321) );
  AO22X1 U3100 ( .A0(n4347), .A1(n1481), .B0(\key_mem[2][56] ), .B1(n4355), 
        .Y(n2065) );
  AO22X1 U3101 ( .A0(n3954), .A1(n1481), .B0(\key_mem[0][56] ), .B1(n3929), 
        .Y(n1809) );
  AO22X1 U3102 ( .A0(n4014), .A1(n1513), .B0(\key_mem[14][88] ), .B1(n4025), 
        .Y(n3569) );
  AO22X1 U3103 ( .A0(n4070), .A1(n1513), .B0(\key_mem[12][88] ), .B1(n4075), 
        .Y(n3313) );
  AO22X1 U3104 ( .A0(n4126), .A1(n1513), .B0(\key_mem[10][88] ), .B1(n4133), 
        .Y(n3057) );
  AO22X1 U3105 ( .A0(n4182), .A1(n1513), .B0(\key_mem[8][88] ), .B1(n4189), 
        .Y(n2801) );
  AO22X1 U3106 ( .A0(n4239), .A1(n1513), .B0(\key_mem[6][88] ), .B1(n4248), 
        .Y(n2545) );
  AO22X1 U3107 ( .A0(n4294), .A1(n1513), .B0(\key_mem[4][88] ), .B1(n4302), 
        .Y(n2289) );
  AO22X1 U3108 ( .A0(n4350), .A1(n1513), .B0(\key_mem[2][88] ), .B1(n4365), 
        .Y(n2033) );
  AO22X1 U3109 ( .A0(n3951), .A1(n1513), .B0(\key_mem[0][88] ), .B1(n3947), 
        .Y(n1777) );
  AO22X1 U3110 ( .A0(n4018), .A1(n1545), .B0(\key_mem[14][120] ), .B1(n4031), 
        .Y(n3537) );
  AO22X1 U3111 ( .A0(n4074), .A1(n1545), .B0(\key_mem[12][120] ), .B1(n4085), 
        .Y(n3281) );
  AO22X1 U3112 ( .A0(n4130), .A1(n1545), .B0(\key_mem[10][120] ), .B1(n4132), 
        .Y(n3025) );
  AO22X1 U3113 ( .A0(n4186), .A1(n1545), .B0(\key_mem[8][120] ), .B1(n4188), 
        .Y(n2769) );
  AO22X1 U3114 ( .A0(n4243), .A1(n1545), .B0(\key_mem[6][120] ), .B1(n4252), 
        .Y(n2513) );
  AO22X1 U3115 ( .A0(n4298), .A1(n1545), .B0(\key_mem[4][120] ), .B1(n4308), 
        .Y(n2257) );
  AO22X1 U3116 ( .A0(n4354), .A1(n1545), .B0(\key_mem[2][120] ), .B1(n4363), 
        .Y(n2001) );
  AO22X1 U3117 ( .A0(n3960), .A1(n1545), .B0(\key_mem[0][120] ), .B1(n3934), 
        .Y(n1745) );
  AO22X1 U3118 ( .A0(n4009), .A1(n1456), .B0(\key_mem[14][31] ), .B1(n4021), 
        .Y(n3626) );
  AO22X1 U3119 ( .A0(n4065), .A1(n1456), .B0(\key_mem[12][31] ), .B1(n4077), 
        .Y(n3370) );
  AO22X1 U3120 ( .A0(n4121), .A1(n1456), .B0(\key_mem[10][31] ), .B1(n4136), 
        .Y(n3114) );
  AO22X1 U3121 ( .A0(n4177), .A1(n1456), .B0(\key_mem[8][31] ), .B1(n4192), 
        .Y(n2858) );
  AO22X1 U3122 ( .A0(n4234), .A1(n1456), .B0(\key_mem[6][31] ), .B1(n4230), 
        .Y(n2602) );
  AO22X1 U3123 ( .A0(n4289), .A1(n1456), .B0(\key_mem[4][31] ), .B1(n4310), 
        .Y(n2346) );
  AO22X1 U3124 ( .A0(n4345), .A1(n1456), .B0(\key_mem[2][31] ), .B1(n4359), 
        .Y(n2090) );
  AO22X1 U3125 ( .A0(n3957), .A1(n1456), .B0(\key_mem[0][31] ), .B1(n1736), 
        .Y(n1834) );
  AO22X1 U3126 ( .A0(n4012), .A1(n1488), .B0(\key_mem[14][63] ), .B1(n4024), 
        .Y(n3594) );
  AO22X1 U3127 ( .A0(n4068), .A1(n1488), .B0(\key_mem[12][63] ), .B1(n4077), 
        .Y(n3338) );
  AO22X1 U3128 ( .A0(n4124), .A1(n1488), .B0(\key_mem[10][63] ), .B1(n4136), 
        .Y(n3082) );
  AO22X1 U3129 ( .A0(n4180), .A1(n1488), .B0(\key_mem[8][63] ), .B1(n4193), 
        .Y(n2826) );
  AO22X1 U3130 ( .A0(n4237), .A1(n1488), .B0(\key_mem[6][63] ), .B1(n4230), 
        .Y(n2570) );
  AO22X1 U3131 ( .A0(n4292), .A1(n1488), .B0(\key_mem[4][63] ), .B1(n4313), 
        .Y(n2314) );
  AO22X1 U3132 ( .A0(n4348), .A1(n1488), .B0(\key_mem[2][63] ), .B1(n4358), 
        .Y(n2058) );
  AO22X1 U3133 ( .A0(n3953), .A1(n1488), .B0(\key_mem[0][63] ), .B1(n3930), 
        .Y(n1802) );
  AO22X1 U3134 ( .A0(n4015), .A1(n1520), .B0(\key_mem[14][95] ), .B1(n4024), 
        .Y(n3562) );
  AO22X1 U3135 ( .A0(n4071), .A1(n1520), .B0(\key_mem[12][95] ), .B1(n4079), 
        .Y(n3306) );
  AO22X1 U3136 ( .A0(n4127), .A1(n1520), .B0(\key_mem[10][95] ), .B1(n4141), 
        .Y(n3050) );
  AO22X1 U3137 ( .A0(n4183), .A1(n1520), .B0(\key_mem[8][95] ), .B1(n4197), 
        .Y(n2794) );
  AO22X1 U3138 ( .A0(n4240), .A1(n1520), .B0(\key_mem[6][95] ), .B1(n4253), 
        .Y(n2538) );
  AO22X1 U3139 ( .A0(n4295), .A1(n1520), .B0(\key_mem[4][95] ), .B1(n4303), 
        .Y(n2282) );
  AO22X1 U3140 ( .A0(n4351), .A1(n1520), .B0(\key_mem[2][95] ), .B1(n4363), 
        .Y(n2026) );
  AO22X1 U3141 ( .A0(n3950), .A1(n1520), .B0(\key_mem[0][95] ), .B1(n3932), 
        .Y(n1770) );
  AO22X1 U3142 ( .A0(n4018), .A1(n1552), .B0(\key_mem[14][127] ), .B1(n4025), 
        .Y(n3530) );
  AO22X1 U3143 ( .A0(n4074), .A1(n1552), .B0(\key_mem[12][127] ), .B1(n4080), 
        .Y(n3274) );
  AO22X1 U3144 ( .A0(n4130), .A1(n1552), .B0(\key_mem[10][127] ), .B1(n4132), 
        .Y(n3018) );
  AO22X1 U3145 ( .A0(n4186), .A1(n1552), .B0(\key_mem[8][127] ), .B1(n4188), 
        .Y(n2762) );
  AO22X1 U3146 ( .A0(n4243), .A1(n1552), .B0(\key_mem[6][127] ), .B1(n730), 
        .Y(n2506) );
  AO22X1 U3147 ( .A0(n4298), .A1(n1552), .B0(\key_mem[4][127] ), .B1(n4300), 
        .Y(n2250) );
  AO22X1 U3148 ( .A0(n4354), .A1(n1552), .B0(\key_mem[2][127] ), .B1(n4358), 
        .Y(n1994) );
  AO22X1 U3149 ( .A0(n3963), .A1(n1552), .B0(\key_mem[0][127] ), .B1(n3930), 
        .Y(n1738) );
  AO22X1 U3150 ( .A0(n4006), .A1(n1426), .B0(\key_mem[14][1] ), .B1(n4019), 
        .Y(n3656) );
  AO22X1 U3151 ( .A0(n4062), .A1(n1426), .B0(\key_mem[12][1] ), .B1(n4075), 
        .Y(n3400) );
  AO22X1 U3152 ( .A0(n4118), .A1(n1426), .B0(\key_mem[10][1] ), .B1(n4131), 
        .Y(n3144) );
  AO22X1 U3153 ( .A0(n4174), .A1(n1426), .B0(\key_mem[8][1] ), .B1(n4187), .Y(
        n2888) );
  AO22X1 U3154 ( .A0(n4231), .A1(n1426), .B0(\key_mem[6][1] ), .B1(n4245), .Y(
        n2632) );
  AO22X1 U3155 ( .A0(n4286), .A1(n1426), .B0(\key_mem[4][1] ), .B1(n4299), .Y(
        n2376) );
  AO22X1 U3156 ( .A0(n4342), .A1(n1426), .B0(\key_mem[2][1] ), .B1(n4355), .Y(
        n2120) );
  AO22X1 U3157 ( .A0(n3960), .A1(n1426), .B0(\key_mem[0][1] ), .B1(n1719), .Y(
        n1864) );
  AO22X1 U3158 ( .A0(n4006), .A1(n1427), .B0(\key_mem[14][2] ), .B1(n4020), 
        .Y(n3655) );
  AO22X1 U3159 ( .A0(n4062), .A1(n1427), .B0(\key_mem[12][2] ), .B1(n4076), 
        .Y(n3399) );
  AO22X1 U3160 ( .A0(n4118), .A1(n1427), .B0(\key_mem[10][2] ), .B1(n4132), 
        .Y(n3143) );
  AO22X1 U3161 ( .A0(n4174), .A1(n1427), .B0(\key_mem[8][2] ), .B1(n4188), .Y(
        n2887) );
  AO22X1 U3162 ( .A0(n4231), .A1(n1427), .B0(\key_mem[6][2] ), .B1(n4246), .Y(
        n2631) );
  AO22X1 U3163 ( .A0(n4286), .A1(n1427), .B0(\key_mem[4][2] ), .B1(n4300), .Y(
        n2375) );
  AO22X1 U3164 ( .A0(n4342), .A1(n1427), .B0(\key_mem[2][2] ), .B1(n4356), .Y(
        n2119) );
  AO22X1 U3165 ( .A0(n3960), .A1(n1427), .B0(\key_mem[0][2] ), .B1(n1719), .Y(
        n1863) );
  AO22X1 U3166 ( .A0(n4006), .A1(n1428), .B0(\key_mem[14][3] ), .B1(n4021), 
        .Y(n3654) );
  AO22X1 U3167 ( .A0(n4062), .A1(n1428), .B0(\key_mem[12][3] ), .B1(n4077), 
        .Y(n3398) );
  AO22X1 U3168 ( .A0(n4118), .A1(n1428), .B0(\key_mem[10][3] ), .B1(n4133), 
        .Y(n3142) );
  AO22X1 U3169 ( .A0(n4174), .A1(n1428), .B0(\key_mem[8][3] ), .B1(n4189), .Y(
        n2886) );
  AO22X1 U3170 ( .A0(n4231), .A1(n1428), .B0(\key_mem[6][3] ), .B1(n4247), .Y(
        n2630) );
  AO22X1 U3171 ( .A0(n4286), .A1(n1428), .B0(\key_mem[4][3] ), .B1(n4301), .Y(
        n2374) );
  AO22X1 U3172 ( .A0(n4342), .A1(n1428), .B0(\key_mem[2][3] ), .B1(n4357), .Y(
        n2118) );
  AO22X1 U3173 ( .A0(n3959), .A1(n1428), .B0(\key_mem[0][3] ), .B1(n1719), .Y(
        n1862) );
  AO22X1 U3174 ( .A0(n4006), .A1(n1429), .B0(\key_mem[14][4] ), .B1(n4022), 
        .Y(n3653) );
  AO22X1 U3175 ( .A0(n4062), .A1(n1429), .B0(\key_mem[12][4] ), .B1(n4078), 
        .Y(n3397) );
  AO22X1 U3176 ( .A0(n4118), .A1(n1429), .B0(\key_mem[10][4] ), .B1(n4134), 
        .Y(n3141) );
  AO22X1 U3177 ( .A0(n4174), .A1(n716), .B0(\key_mem[8][4] ), .B1(n4190), .Y(
        n2885) );
  AO22X1 U3178 ( .A0(n4231), .A1(n716), .B0(\key_mem[6][4] ), .B1(n4248), .Y(
        n2629) );
  AO22X1 U3179 ( .A0(n4286), .A1(n716), .B0(\key_mem[4][4] ), .B1(n4302), .Y(
        n2373) );
  AO22X1 U3180 ( .A0(n4342), .A1(n716), .B0(\key_mem[2][4] ), .B1(n4358), .Y(
        n2117) );
  AO22X1 U3181 ( .A0(n3959), .A1(n716), .B0(\key_mem[0][4] ), .B1(n1719), .Y(
        n1861) );
  AO22X1 U3182 ( .A0(n4006), .A1(n1430), .B0(\key_mem[14][5] ), .B1(n4023), 
        .Y(n3652) );
  AO22X1 U3183 ( .A0(n4062), .A1(n1430), .B0(\key_mem[12][5] ), .B1(n4079), 
        .Y(n3396) );
  AO22X1 U3184 ( .A0(n4118), .A1(n1430), .B0(\key_mem[10][5] ), .B1(n4135), 
        .Y(n3140) );
  AO22X1 U3185 ( .A0(n4174), .A1(n1430), .B0(\key_mem[8][5] ), .B1(n4191), .Y(
        n2884) );
  AO22X1 U3186 ( .A0(n4231), .A1(n1430), .B0(\key_mem[6][5] ), .B1(n4249), .Y(
        n2628) );
  AO22X1 U3187 ( .A0(n4286), .A1(n1430), .B0(\key_mem[4][5] ), .B1(n4303), .Y(
        n2372) );
  AO22X1 U3188 ( .A0(n4342), .A1(n1430), .B0(\key_mem[2][5] ), .B1(n4359), .Y(
        n2116) );
  AO22X1 U3189 ( .A0(n3959), .A1(n1430), .B0(\key_mem[0][5] ), .B1(n1719), .Y(
        n1860) );
  AO22X1 U3190 ( .A0(n4006), .A1(n1432), .B0(\key_mem[14][7] ), .B1(n4025), 
        .Y(n3650) );
  AO22X1 U3191 ( .A0(n4062), .A1(n1432), .B0(\key_mem[12][7] ), .B1(n4081), 
        .Y(n3394) );
  AO22X1 U3192 ( .A0(n4118), .A1(n1432), .B0(\key_mem[10][7] ), .B1(n4137), 
        .Y(n3138) );
  AO22X1 U3193 ( .A0(n4174), .A1(n1432), .B0(\key_mem[8][7] ), .B1(n4193), .Y(
        n2882) );
  AO22X1 U3194 ( .A0(n4231), .A1(n1432), .B0(\key_mem[6][7] ), .B1(n4251), .Y(
        n2626) );
  AO22X1 U3195 ( .A0(n4286), .A1(n1432), .B0(\key_mem[4][7] ), .B1(n4305), .Y(
        n2370) );
  AO22X1 U3196 ( .A0(n4342), .A1(n1432), .B0(\key_mem[2][7] ), .B1(n4361), .Y(
        n2114) );
  AO22X1 U3197 ( .A0(n3959), .A1(n1432), .B0(\key_mem[0][7] ), .B1(n1719), .Y(
        n1858) );
  AO22X1 U3198 ( .A0(n4007), .A1(n1435), .B0(\key_mem[14][10] ), .B1(n4027), 
        .Y(n3647) );
  AO22X1 U3199 ( .A0(n4063), .A1(n1435), .B0(\key_mem[12][10] ), .B1(n738), 
        .Y(n3391) );
  AO22X1 U3200 ( .A0(n4119), .A1(n1435), .B0(\key_mem[10][10] ), .B1(n4140), 
        .Y(n3135) );
  AO22X1 U3201 ( .A0(n4175), .A1(n1435), .B0(\key_mem[8][10] ), .B1(n4196), 
        .Y(n2879) );
  AO22X1 U3202 ( .A0(n4232), .A1(n1435), .B0(\key_mem[6][10] ), .B1(n4251), 
        .Y(n2623) );
  AO22X1 U3203 ( .A0(n4287), .A1(n1435), .B0(\key_mem[4][10] ), .B1(n4308), 
        .Y(n2367) );
  AO22X1 U3204 ( .A0(n4343), .A1(n1435), .B0(\key_mem[2][10] ), .B1(n4364), 
        .Y(n2111) );
  AO22X1 U3205 ( .A0(n3959), .A1(n1435), .B0(\key_mem[0][10] ), .B1(n1719), 
        .Y(n1855) );
  AO22X1 U3206 ( .A0(n4007), .A1(n1438), .B0(\key_mem[14][13] ), .B1(n4032), 
        .Y(n3644) );
  AO22X1 U3207 ( .A0(n4063), .A1(n1438), .B0(\key_mem[12][13] ), .B1(n4087), 
        .Y(n3388) );
  AO22X1 U3208 ( .A0(n4119), .A1(n1438), .B0(\key_mem[10][13] ), .B1(n4144), 
        .Y(n3132) );
  AO22X1 U3209 ( .A0(n4175), .A1(n1438), .B0(\key_mem[8][13] ), .B1(n4200), 
        .Y(n2876) );
  AO22X1 U3210 ( .A0(n4232), .A1(n1438), .B0(\key_mem[6][13] ), .B1(n730), .Y(
        n2620) );
  AO22X1 U3211 ( .A0(n4287), .A1(n1438), .B0(\key_mem[4][13] ), .B1(n4307), 
        .Y(n2364) );
  AO22X1 U3212 ( .A0(n4343), .A1(n1438), .B0(\key_mem[2][13] ), .B1(n4356), 
        .Y(n2108) );
  AO22X1 U3213 ( .A0(n3958), .A1(n1438), .B0(\key_mem[0][13] ), .B1(n1720), 
        .Y(n1852) );
  AO22X1 U3214 ( .A0(n4007), .A1(n1443), .B0(\key_mem[14][18] ), .B1(n4033), 
        .Y(n3639) );
  AO22X1 U3215 ( .A0(n4063), .A1(n1443), .B0(\key_mem[12][18] ), .B1(n4088), 
        .Y(n3383) );
  AO22X1 U3216 ( .A0(n4119), .A1(n1443), .B0(\key_mem[10][18] ), .B1(n4145), 
        .Y(n3127) );
  AO22X1 U3217 ( .A0(n4175), .A1(n1443), .B0(\key_mem[8][18] ), .B1(n4201), 
        .Y(n2871) );
  AO22X1 U3218 ( .A0(n4232), .A1(n1443), .B0(\key_mem[6][18] ), .B1(n730), .Y(
        n2615) );
  AO22X1 U3219 ( .A0(n4287), .A1(n1443), .B0(\key_mem[4][18] ), .B1(n4311), 
        .Y(n2359) );
  AO22X1 U3220 ( .A0(n4343), .A1(n1443), .B0(\key_mem[2][18] ), .B1(n4355), 
        .Y(n2103) );
  AO22X1 U3221 ( .A0(n3958), .A1(n1443), .B0(\key_mem[0][18] ), .B1(n1720), 
        .Y(n1847) );
  AO22X1 U3222 ( .A0(n4008), .A1(n1447), .B0(\key_mem[14][22] ), .B1(n4026), 
        .Y(n3635) );
  AO22X1 U3223 ( .A0(n4064), .A1(n1447), .B0(\key_mem[12][22] ), .B1(n4089), 
        .Y(n3379) );
  AO22X1 U3224 ( .A0(n4120), .A1(n1447), .B0(\key_mem[10][22] ), .B1(n4143), 
        .Y(n3123) );
  AO22X1 U3225 ( .A0(n4176), .A1(n1447), .B0(\key_mem[8][22] ), .B1(n4199), 
        .Y(n2867) );
  AO22X1 U3226 ( .A0(n4233), .A1(n1447), .B0(\key_mem[6][22] ), .B1(n4250), 
        .Y(n2611) );
  AO22X1 U3227 ( .A0(n4288), .A1(n1447), .B0(\key_mem[4][22] ), .B1(n4312), 
        .Y(n2355) );
  AO22X1 U3228 ( .A0(n4344), .A1(n1447), .B0(\key_mem[2][22] ), .B1(n4358), 
        .Y(n2099) );
  AO22X1 U3229 ( .A0(n3958), .A1(n1447), .B0(\key_mem[0][22] ), .B1(n1728), 
        .Y(n1843) );
  AO22X1 U3230 ( .A0(n4009), .A1(n1458), .B0(\key_mem[14][33] ), .B1(n4020), 
        .Y(n3624) );
  AO22X1 U3231 ( .A0(n4065), .A1(n1458), .B0(\key_mem[12][33] ), .B1(n4089), 
        .Y(n3368) );
  AO22X1 U3232 ( .A0(n4121), .A1(n1458), .B0(\key_mem[10][33] ), .B1(n4137), 
        .Y(n3112) );
  AO22X1 U3233 ( .A0(n4177), .A1(n1458), .B0(\key_mem[8][33] ), .B1(n4193), 
        .Y(n2856) );
  AO22X1 U3234 ( .A0(n4234), .A1(n1458), .B0(\key_mem[6][33] ), .B1(n4255), 
        .Y(n2600) );
  AO22X1 U3235 ( .A0(n4289), .A1(n1458), .B0(\key_mem[4][33] ), .B1(n4304), 
        .Y(n2344) );
  AO22X1 U3236 ( .A0(n4345), .A1(n1458), .B0(\key_mem[2][33] ), .B1(n4358), 
        .Y(n2088) );
  AO22X1 U3237 ( .A0(n3956), .A1(n1458), .B0(\key_mem[0][33] ), .B1(n1736), 
        .Y(n1832) );
  AO22X1 U3238 ( .A0(n4009), .A1(n1459), .B0(\key_mem[14][34] ), .B1(n4031), 
        .Y(n3623) );
  AO22X1 U3239 ( .A0(n4065), .A1(n1459), .B0(\key_mem[12][34] ), .B1(n4081), 
        .Y(n3367) );
  AO22X1 U3240 ( .A0(n4121), .A1(n1459), .B0(\key_mem[10][34] ), .B1(n4143), 
        .Y(n3111) );
  AO22X1 U3241 ( .A0(n4177), .A1(n1459), .B0(\key_mem[8][34] ), .B1(n4199), 
        .Y(n2855) );
  AO22X1 U3242 ( .A0(n4234), .A1(n1459), .B0(\key_mem[6][34] ), .B1(n4256), 
        .Y(n2599) );
  AO22X1 U3243 ( .A0(n4289), .A1(n1459), .B0(\key_mem[4][34] ), .B1(n4306), 
        .Y(n2343) );
  AO22X1 U3244 ( .A0(n4345), .A1(n1459), .B0(\key_mem[2][34] ), .B1(n4367), 
        .Y(n2087) );
  AO22X1 U3245 ( .A0(n3956), .A1(n1459), .B0(\key_mem[0][34] ), .B1(n1736), 
        .Y(n1831) );
  AO22X1 U3246 ( .A0(n4009), .A1(n1460), .B0(\key_mem[14][35] ), .B1(n4020), 
        .Y(n3622) );
  AO22X1 U3247 ( .A0(n4065), .A1(n1460), .B0(\key_mem[12][35] ), .B1(n4076), 
        .Y(n3366) );
  AO22X1 U3248 ( .A0(n4121), .A1(n1460), .B0(\key_mem[10][35] ), .B1(n4144), 
        .Y(n3110) );
  AO22X1 U3249 ( .A0(n4177), .A1(n1460), .B0(\key_mem[8][35] ), .B1(n4200), 
        .Y(n2854) );
  AO22X1 U3250 ( .A0(n4234), .A1(n1460), .B0(\key_mem[6][35] ), .B1(n4255), 
        .Y(n2598) );
  AO22X1 U3251 ( .A0(n4289), .A1(n1460), .B0(\key_mem[4][35] ), .B1(n4306), 
        .Y(n2342) );
  AO22X1 U3252 ( .A0(n4345), .A1(n1460), .B0(\key_mem[2][35] ), .B1(n4368), 
        .Y(n2086) );
  AO22X1 U3253 ( .A0(n3956), .A1(n1460), .B0(\key_mem[0][35] ), .B1(n1736), 
        .Y(n1830) );
  AO22X1 U3254 ( .A0(n4009), .A1(n1461), .B0(\key_mem[14][36] ), .B1(n4032), 
        .Y(n3621) );
  AO22X1 U3255 ( .A0(n4065), .A1(n1461), .B0(\key_mem[12][36] ), .B1(n4087), 
        .Y(n3365) );
  AO22X1 U3256 ( .A0(n4121), .A1(n1461), .B0(\key_mem[10][36] ), .B1(n4145), 
        .Y(n3109) );
  AO22X1 U3257 ( .A0(n4177), .A1(n1461), .B0(\key_mem[8][36] ), .B1(n4201), 
        .Y(n2853) );
  AO22X1 U3258 ( .A0(n4234), .A1(n1461), .B0(\key_mem[6][36] ), .B1(n4255), 
        .Y(n2597) );
  AO22X1 U3259 ( .A0(n4289), .A1(n1461), .B0(\key_mem[4][36] ), .B1(n4305), 
        .Y(n2341) );
  AO22X1 U3260 ( .A0(n4345), .A1(n1461), .B0(\key_mem[2][36] ), .B1(n4369), 
        .Y(n2085) );
  AO22X1 U3261 ( .A0(n3956), .A1(n1461), .B0(\key_mem[0][36] ), .B1(n1736), 
        .Y(n1829) );
  AO22X1 U3262 ( .A0(n4009), .A1(n1462), .B0(\key_mem[14][37] ), .B1(n4019), 
        .Y(n3620) );
  AO22X1 U3263 ( .A0(n4065), .A1(n1462), .B0(\key_mem[12][37] ), .B1(n4076), 
        .Y(n3364) );
  AO22X1 U3264 ( .A0(n4121), .A1(n1462), .B0(\key_mem[10][37] ), .B1(n4144), 
        .Y(n3108) );
  AO22X1 U3265 ( .A0(n4177), .A1(n1462), .B0(\key_mem[8][37] ), .B1(n4200), 
        .Y(n2852) );
  AO22X1 U3266 ( .A0(n4234), .A1(n1462), .B0(\key_mem[6][37] ), .B1(n4256), 
        .Y(n2596) );
  AO22X1 U3267 ( .A0(n4289), .A1(n1462), .B0(\key_mem[4][37] ), .B1(n4307), 
        .Y(n2340) );
  AO22X1 U3268 ( .A0(n4345), .A1(n1462), .B0(\key_mem[2][37] ), .B1(n4357), 
        .Y(n2084) );
  AO22X1 U3269 ( .A0(n3956), .A1(n1462), .B0(\key_mem[0][37] ), .B1(n1736), 
        .Y(n1828) );
  AO22X1 U3270 ( .A0(n4009), .A1(n1464), .B0(\key_mem[14][39] ), .B1(n4033), 
        .Y(n3618) );
  AO22X1 U3271 ( .A0(n4065), .A1(n1464), .B0(\key_mem[12][39] ), .B1(n4086), 
        .Y(n3362) );
  AO22X1 U3272 ( .A0(n4121), .A1(n1464), .B0(\key_mem[10][39] ), .B1(n4144), 
        .Y(n3106) );
  AO22X1 U3273 ( .A0(n4177), .A1(n1464), .B0(\key_mem[8][39] ), .B1(n4200), 
        .Y(n2850) );
  AO22X1 U3274 ( .A0(n4234), .A1(n1464), .B0(\key_mem[6][39] ), .B1(n4244), 
        .Y(n2594) );
  AO22X1 U3275 ( .A0(n4289), .A1(n1464), .B0(\key_mem[4][39] ), .B1(n4302), 
        .Y(n2338) );
  AO22X1 U3276 ( .A0(n4345), .A1(n1464), .B0(\key_mem[2][39] ), .B1(n4367), 
        .Y(n2082) );
  AO22X1 U3277 ( .A0(n3956), .A1(n1464), .B0(\key_mem[0][39] ), .B1(n1736), 
        .Y(n1826) );
  AO22X1 U3278 ( .A0(n4010), .A1(n1467), .B0(\key_mem[14][42] ), .B1(n4033), 
        .Y(n3615) );
  AO22X1 U3279 ( .A0(n4066), .A1(n1467), .B0(\key_mem[12][42] ), .B1(n4083), 
        .Y(n3359) );
  AO22X1 U3280 ( .A0(n4122), .A1(n1467), .B0(\key_mem[10][42] ), .B1(n4135), 
        .Y(n3103) );
  AO22X1 U3281 ( .A0(n4178), .A1(n1467), .B0(\key_mem[8][42] ), .B1(n4191), 
        .Y(n2847) );
  AO22X1 U3282 ( .A0(n4235), .A1(n1467), .B0(\key_mem[6][42] ), .B1(n4244), 
        .Y(n2591) );
  AO22X1 U3283 ( .A0(n4290), .A1(n1467), .B0(\key_mem[4][42] ), .B1(n4305), 
        .Y(n2335) );
  AO22X1 U3284 ( .A0(n4346), .A1(n1467), .B0(\key_mem[2][42] ), .B1(n4368), 
        .Y(n2079) );
  AO22X1 U3285 ( .A0(n3956), .A1(n1467), .B0(\key_mem[0][42] ), .B1(n3928), 
        .Y(n1823) );
  AO22X1 U3286 ( .A0(n4010), .A1(n1470), .B0(\key_mem[14][45] ), .B1(n4033), 
        .Y(n3612) );
  AO22X1 U3287 ( .A0(n4066), .A1(n1470), .B0(\key_mem[12][45] ), .B1(n4082), 
        .Y(n3356) );
  AO22X1 U3288 ( .A0(n4122), .A1(n1470), .B0(\key_mem[10][45] ), .B1(n4142), 
        .Y(n3100) );
  AO22X1 U3289 ( .A0(n4178), .A1(n1470), .B0(\key_mem[8][45] ), .B1(n4198), 
        .Y(n2844) );
  AO22X1 U3290 ( .A0(n4235), .A1(n1470), .B0(\key_mem[6][45] ), .B1(n4257), 
        .Y(n2588) );
  AO22X1 U3291 ( .A0(n4290), .A1(n1470), .B0(\key_mem[4][45] ), .B1(n4312), 
        .Y(n2332) );
  AO22X1 U3292 ( .A0(n4346), .A1(n1470), .B0(\key_mem[2][45] ), .B1(n4369), 
        .Y(n2076) );
  AO22X1 U3293 ( .A0(n3955), .A1(n1470), .B0(\key_mem[0][45] ), .B1(n3928), 
        .Y(n1820) );
  AO22X1 U3294 ( .A0(n4011), .A1(n1475), .B0(\key_mem[14][50] ), .B1(n4031), 
        .Y(n3607) );
  AO22X1 U3295 ( .A0(n4067), .A1(n1475), .B0(\key_mem[12][50] ), .B1(n4086), 
        .Y(n3351) );
  AO22X1 U3296 ( .A0(n4123), .A1(n1475), .B0(\key_mem[10][50] ), .B1(n4134), 
        .Y(n3095) );
  AO22X1 U3297 ( .A0(n4179), .A1(n1475), .B0(\key_mem[8][50] ), .B1(n4190), 
        .Y(n2839) );
  AO22X1 U3298 ( .A0(n4236), .A1(n1475), .B0(\key_mem[6][50] ), .B1(n4257), 
        .Y(n2583) );
  AO22X1 U3299 ( .A0(n4291), .A1(n1475), .B0(\key_mem[4][50] ), .B1(n4313), 
        .Y(n2327) );
  AO22X1 U3300 ( .A0(n4347), .A1(n1475), .B0(\key_mem[2][50] ), .B1(n4357), 
        .Y(n2071) );
  AO22X1 U3301 ( .A0(n3955), .A1(n1475), .B0(\key_mem[0][50] ), .B1(n3928), 
        .Y(n1815) );
  AO22X1 U3302 ( .A0(n4011), .A1(n1478), .B0(\key_mem[14][53] ), .B1(n4025), 
        .Y(n3604) );
  AO22X1 U3303 ( .A0(n4067), .A1(n1478), .B0(\key_mem[12][53] ), .B1(n4076), 
        .Y(n3348) );
  AO22X1 U3304 ( .A0(n4123), .A1(n1478), .B0(\key_mem[10][53] ), .B1(n4134), 
        .Y(n3092) );
  AO22X1 U3305 ( .A0(n4179), .A1(n1478), .B0(\key_mem[8][53] ), .B1(n4190), 
        .Y(n2836) );
  AO22X1 U3306 ( .A0(n4236), .A1(n1478), .B0(\key_mem[6][53] ), .B1(n4250), 
        .Y(n2580) );
  AO22X1 U3307 ( .A0(n4291), .A1(n1478), .B0(\key_mem[4][53] ), .B1(n4300), 
        .Y(n2324) );
  AO22X1 U3308 ( .A0(n4347), .A1(n1478), .B0(\key_mem[2][53] ), .B1(n4359), 
        .Y(n2068) );
  AO22X1 U3309 ( .A0(n3954), .A1(n1478), .B0(\key_mem[0][53] ), .B1(n3929), 
        .Y(n1812) );
  AO22X1 U3310 ( .A0(n4011), .A1(n1480), .B0(\key_mem[14][55] ), .B1(n4023), 
        .Y(n3602) );
  AO22X1 U3311 ( .A0(n4067), .A1(n1480), .B0(\key_mem[12][55] ), .B1(n4075), 
        .Y(n3346) );
  AO22X1 U3312 ( .A0(n4123), .A1(n1480), .B0(\key_mem[10][55] ), .B1(n4136), 
        .Y(n3090) );
  AO22X1 U3313 ( .A0(n4179), .A1(n1480), .B0(\key_mem[8][55] ), .B1(n4192), 
        .Y(n2834) );
  AO22X1 U3314 ( .A0(n4236), .A1(n1480), .B0(\key_mem[6][55] ), .B1(n4249), 
        .Y(n2578) );
  AO22X1 U3315 ( .A0(n4291), .A1(n1480), .B0(\key_mem[4][55] ), .B1(n4303), 
        .Y(n2322) );
  AO22X1 U3316 ( .A0(n4347), .A1(n1480), .B0(\key_mem[2][55] ), .B1(n722), .Y(
        n2066) );
  AO22X1 U3317 ( .A0(n3954), .A1(n1480), .B0(\key_mem[0][55] ), .B1(n3929), 
        .Y(n1810) );
  AO22X1 U3318 ( .A0(n4012), .A1(n1490), .B0(\key_mem[14][65] ), .B1(n4022), 
        .Y(n3592) );
  AO22X1 U3319 ( .A0(n4068), .A1(n1490), .B0(\key_mem[12][65] ), .B1(n4076), 
        .Y(n3336) );
  AO22X1 U3320 ( .A0(n4124), .A1(n1490), .B0(\key_mem[10][65] ), .B1(n4135), 
        .Y(n3080) );
  AO22X1 U3321 ( .A0(n4180), .A1(n1490), .B0(\key_mem[8][65] ), .B1(n4192), 
        .Y(n2824) );
  AO22X1 U3322 ( .A0(n4237), .A1(n1490), .B0(\key_mem[6][65] ), .B1(n4244), 
        .Y(n2568) );
  AO22X1 U3323 ( .A0(n4292), .A1(n1490), .B0(\key_mem[4][65] ), .B1(n4306), 
        .Y(n2312) );
  AO22X1 U3324 ( .A0(n4348), .A1(n1490), .B0(\key_mem[2][65] ), .B1(n4363), 
        .Y(n2056) );
  AO22X1 U3325 ( .A0(n3953), .A1(n1490), .B0(\key_mem[0][65] ), .B1(n3930), 
        .Y(n1800) );
  AO22X1 U3326 ( .A0(n4012), .A1(n1491), .B0(\key_mem[14][66] ), .B1(n4021), 
        .Y(n3591) );
  AO22X1 U3327 ( .A0(n4068), .A1(n1491), .B0(\key_mem[12][66] ), .B1(n4075), 
        .Y(n3335) );
  AO22X1 U3328 ( .A0(n4124), .A1(n1491), .B0(\key_mem[10][66] ), .B1(n4134), 
        .Y(n3079) );
  AO22X1 U3329 ( .A0(n4180), .A1(n1491), .B0(\key_mem[8][66] ), .B1(n4191), 
        .Y(n2823) );
  AO22X1 U3330 ( .A0(n4237), .A1(n1491), .B0(\key_mem[6][66] ), .B1(n730), .Y(
        n2567) );
  AO22X1 U3331 ( .A0(n4292), .A1(n1491), .B0(\key_mem[4][66] ), .B1(n4311), 
        .Y(n2311) );
  AO22X1 U3332 ( .A0(n4348), .A1(n1491), .B0(\key_mem[2][66] ), .B1(n722), .Y(
        n2055) );
  AO22X1 U3333 ( .A0(n3953), .A1(n1491), .B0(\key_mem[0][66] ), .B1(n3930), 
        .Y(n1799) );
  AO22X1 U3334 ( .A0(n4012), .A1(n1492), .B0(\key_mem[14][67] ), .B1(n4025), 
        .Y(n3590) );
  AO22X1 U3335 ( .A0(n4068), .A1(n1492), .B0(\key_mem[12][67] ), .B1(n4083), 
        .Y(n3334) );
  AO22X1 U3336 ( .A0(n4124), .A1(n1492), .B0(\key_mem[10][67] ), .B1(n4133), 
        .Y(n3078) );
  AO22X1 U3337 ( .A0(n4180), .A1(n1492), .B0(\key_mem[8][67] ), .B1(n4190), 
        .Y(n2822) );
  AO22X1 U3338 ( .A0(n4237), .A1(n1492), .B0(\key_mem[6][67] ), .B1(n730), .Y(
        n2566) );
  AO22X1 U3339 ( .A0(n4292), .A1(n1492), .B0(\key_mem[4][67] ), .B1(n4312), 
        .Y(n2310) );
  AO22X1 U3340 ( .A0(n4348), .A1(n1492), .B0(\key_mem[2][67] ), .B1(n4367), 
        .Y(n2054) );
  AO22X1 U3341 ( .A0(n3953), .A1(n1492), .B0(\key_mem[0][67] ), .B1(n3930), 
        .Y(n1798) );
  AO22X1 U3342 ( .A0(n4012), .A1(n1493), .B0(\key_mem[14][68] ), .B1(n4028), 
        .Y(n3589) );
  AO22X1 U3343 ( .A0(n4068), .A1(n1493), .B0(\key_mem[12][68] ), .B1(n4082), 
        .Y(n3333) );
  AO22X1 U3344 ( .A0(n4124), .A1(n1493), .B0(\key_mem[10][68] ), .B1(n4131), 
        .Y(n3077) );
  AO22X1 U3345 ( .A0(n4180), .A1(n1493), .B0(\key_mem[8][68] ), .B1(n4189), 
        .Y(n2821) );
  AO22X1 U3346 ( .A0(n4237), .A1(n1493), .B0(\key_mem[6][68] ), .B1(n730), .Y(
        n2565) );
  AO22X1 U3347 ( .A0(n4292), .A1(n1493), .B0(\key_mem[4][68] ), .B1(n4313), 
        .Y(n2309) );
  AO22X1 U3348 ( .A0(n4348), .A1(n1493), .B0(\key_mem[2][68] ), .B1(n4368), 
        .Y(n2053) );
  AO22X1 U3349 ( .A0(n3953), .A1(n1493), .B0(\key_mem[0][68] ), .B1(n3930), 
        .Y(n1797) );
  AO22X1 U3350 ( .A0(n4012), .A1(n1494), .B0(\key_mem[14][69] ), .B1(n4027), 
        .Y(n3588) );
  AO22X1 U3351 ( .A0(n4068), .A1(n1494), .B0(\key_mem[12][69] ), .B1(n4081), 
        .Y(n3332) );
  AO22X1 U3352 ( .A0(n4124), .A1(n1494), .B0(\key_mem[10][69] ), .B1(n4132), 
        .Y(n3076) );
  AO22X1 U3353 ( .A0(n4180), .A1(n1494), .B0(\key_mem[8][69] ), .B1(n4187), 
        .Y(n2820) );
  AO22X1 U3354 ( .A0(n4237), .A1(n1494), .B0(\key_mem[6][69] ), .B1(n4250), 
        .Y(n2564) );
  AO22X1 U3355 ( .A0(n4292), .A1(n1494), .B0(\key_mem[4][69] ), .B1(n4310), 
        .Y(n2308) );
  AO22X1 U3356 ( .A0(n4348), .A1(n1494), .B0(\key_mem[2][69] ), .B1(n4369), 
        .Y(n2052) );
  AO22X1 U3357 ( .A0(n3953), .A1(n1494), .B0(\key_mem[0][69] ), .B1(n3931), 
        .Y(n1796) );
  AO22X1 U3358 ( .A0(n4013), .A1(n1496), .B0(\key_mem[14][71] ), .B1(n4029), 
        .Y(n3586) );
  AO22X1 U3359 ( .A0(n4069), .A1(n1496), .B0(\key_mem[12][71] ), .B1(n4081), 
        .Y(n3330) );
  AO22X1 U3360 ( .A0(n4125), .A1(n1496), .B0(\key_mem[10][71] ), .B1(n4139), 
        .Y(n3074) );
  AO22X1 U3361 ( .A0(n4181), .A1(n1496), .B0(\key_mem[8][71] ), .B1(n4188), 
        .Y(n2818) );
  AO22X1 U3362 ( .A0(n4238), .A1(n1496), .B0(\key_mem[6][71] ), .B1(n4249), 
        .Y(n2562) );
  AO22X1 U3363 ( .A0(n4293), .A1(n1496), .B0(\key_mem[4][71] ), .B1(n4307), 
        .Y(n2306) );
  AO22X1 U3364 ( .A0(n4349), .A1(n1496), .B0(\key_mem[2][71] ), .B1(n4362), 
        .Y(n2050) );
  AO22X1 U3365 ( .A0(n3953), .A1(n1496), .B0(\key_mem[0][71] ), .B1(n3931), 
        .Y(n1794) );
  AO22X1 U3366 ( .A0(n4013), .A1(n1499), .B0(\key_mem[14][74] ), .B1(n4019), 
        .Y(n3583) );
  AO22X1 U3367 ( .A0(n4069), .A1(n1499), .B0(\key_mem[12][74] ), .B1(n4082), 
        .Y(n3327) );
  AO22X1 U3368 ( .A0(n4125), .A1(n1499), .B0(\key_mem[10][74] ), .B1(n4132), 
        .Y(n3071) );
  AO22X1 U3369 ( .A0(n4181), .A1(n1499), .B0(\key_mem[8][74] ), .B1(n4188), 
        .Y(n2815) );
  AO22X1 U3370 ( .A0(n4238), .A1(n1499), .B0(\key_mem[6][74] ), .B1(n4249), 
        .Y(n2559) );
  AO22X1 U3371 ( .A0(n4293), .A1(n1499), .B0(\key_mem[4][74] ), .B1(n4307), 
        .Y(n2303) );
  AO22X1 U3372 ( .A0(n4349), .A1(n1499), .B0(\key_mem[2][74] ), .B1(n4366), 
        .Y(n2047) );
  AO22X1 U3373 ( .A0(n3952), .A1(n1499), .B0(\key_mem[0][74] ), .B1(n3931), 
        .Y(n1791) );
  AO22X1 U3374 ( .A0(n4013), .A1(n1502), .B0(\key_mem[14][77] ), .B1(n4028), 
        .Y(n3580) );
  AO22X1 U3375 ( .A0(n4069), .A1(n1502), .B0(\key_mem[12][77] ), .B1(n4081), 
        .Y(n3324) );
  AO22X1 U3376 ( .A0(n4125), .A1(n1502), .B0(\key_mem[10][77] ), .B1(n4139), 
        .Y(n3068) );
  AO22X1 U3377 ( .A0(n4181), .A1(n1502), .B0(\key_mem[8][77] ), .B1(n4195), 
        .Y(n2812) );
  AO22X1 U3378 ( .A0(n4238), .A1(n1502), .B0(\key_mem[6][77] ), .B1(n4247), 
        .Y(n2556) );
  AO22X1 U3379 ( .A0(n4293), .A1(n1502), .B0(\key_mem[4][77] ), .B1(n4305), 
        .Y(n2300) );
  AO22X1 U3380 ( .A0(n4349), .A1(n1502), .B0(\key_mem[2][77] ), .B1(n4366), 
        .Y(n2044) );
  AO22X1 U3381 ( .A0(n3952), .A1(n1502), .B0(\key_mem[0][77] ), .B1(n3931), 
        .Y(n1788) );
  AO22X1 U3382 ( .A0(n4013), .A1(n1504), .B0(\key_mem[14][79] ), .B1(n4027), 
        .Y(n3578) );
  AO22X1 U3383 ( .A0(n4069), .A1(n1504), .B0(\key_mem[12][79] ), .B1(n4083), 
        .Y(n3322) );
  AO22X1 U3384 ( .A0(n4125), .A1(n1504), .B0(\key_mem[10][79] ), .B1(n4138), 
        .Y(n3066) );
  AO22X1 U3385 ( .A0(n4181), .A1(n1504), .B0(\key_mem[8][79] ), .B1(n4194), 
        .Y(n2810) );
  AO22X1 U3386 ( .A0(n4238), .A1(n1504), .B0(\key_mem[6][79] ), .B1(n4246), 
        .Y(n2554) );
  AO22X1 U3387 ( .A0(n4293), .A1(n1504), .B0(\key_mem[4][79] ), .B1(n4303), 
        .Y(n2298) );
  AO22X1 U3388 ( .A0(n4349), .A1(n1504), .B0(\key_mem[2][79] ), .B1(n4366), 
        .Y(n2042) );
  AO22X1 U3389 ( .A0(n3952), .A1(n1504), .B0(\key_mem[0][79] ), .B1(n1717), 
        .Y(n1786) );
  AO22X1 U3390 ( .A0(n4014), .A1(n1506), .B0(\key_mem[14][81] ), .B1(n4029), 
        .Y(n3576) );
  AO22X1 U3391 ( .A0(n4070), .A1(n1506), .B0(\key_mem[12][81] ), .B1(n4075), 
        .Y(n3320) );
  AO22X1 U3392 ( .A0(n4126), .A1(n1506), .B0(\key_mem[10][81] ), .B1(n4137), 
        .Y(n3064) );
  AO22X1 U3393 ( .A0(n4182), .A1(n1506), .B0(\key_mem[8][81] ), .B1(n4193), 
        .Y(n2808) );
  AO22X1 U3394 ( .A0(n4239), .A1(n1506), .B0(\key_mem[6][81] ), .B1(n4248), 
        .Y(n2552) );
  AO22X1 U3395 ( .A0(n4294), .A1(n1506), .B0(\key_mem[4][81] ), .B1(n4302), 
        .Y(n2296) );
  AO22X1 U3396 ( .A0(n4350), .A1(n1506), .B0(\key_mem[2][81] ), .B1(n4366), 
        .Y(n2040) );
  AO22X1 U3397 ( .A0(n3952), .A1(n1506), .B0(\key_mem[0][81] ), .B1(n5761), 
        .Y(n1784) );
  AO22X1 U3398 ( .A0(n4014), .A1(n1507), .B0(\key_mem[14][82] ), .B1(n4020), 
        .Y(n3575) );
  AO22X1 U3399 ( .A0(n4070), .A1(n1507), .B0(\key_mem[12][82] ), .B1(n4079), 
        .Y(n3319) );
  AO22X1 U3400 ( .A0(n4126), .A1(n1507), .B0(\key_mem[10][82] ), .B1(n4136), 
        .Y(n3063) );
  AO22X1 U3401 ( .A0(n4182), .A1(n1507), .B0(\key_mem[8][82] ), .B1(n4190), 
        .Y(n2807) );
  AO22X1 U3402 ( .A0(n4239), .A1(n1507), .B0(\key_mem[6][82] ), .B1(n4249), 
        .Y(n2551) );
  AO22X1 U3403 ( .A0(n4294), .A1(n1507), .B0(\key_mem[4][82] ), .B1(n4301), 
        .Y(n2295) );
  AO22X1 U3404 ( .A0(n4350), .A1(n1507), .B0(\key_mem[2][82] ), .B1(n4366), 
        .Y(n2039) );
  AO22X1 U3405 ( .A0(n3952), .A1(n1507), .B0(\key_mem[0][82] ), .B1(n5761), 
        .Y(n1783) );
  AO22X1 U3406 ( .A0(n4014), .A1(n1509), .B0(\key_mem[14][84] ), .B1(n4023), 
        .Y(n3573) );
  AO22X1 U3407 ( .A0(n4070), .A1(n1509), .B0(\key_mem[12][84] ), .B1(n4080), 
        .Y(n3317) );
  AO22X1 U3408 ( .A0(n4126), .A1(n1509), .B0(\key_mem[10][84] ), .B1(n4132), 
        .Y(n3061) );
  AO22X1 U3409 ( .A0(n4182), .A1(n1509), .B0(\key_mem[8][84] ), .B1(n4188), 
        .Y(n2805) );
  AO22X1 U3410 ( .A0(n4239), .A1(n1509), .B0(\key_mem[6][84] ), .B1(n4245), 
        .Y(n2549) );
  AO22X1 U3411 ( .A0(n4294), .A1(n1509), .B0(\key_mem[4][84] ), .B1(n4301), 
        .Y(n2293) );
  AO22X1 U3412 ( .A0(n4350), .A1(n1509), .B0(\key_mem[2][84] ), .B1(n4364), 
        .Y(n2037) );
  AO22X1 U3413 ( .A0(n3951), .A1(n1509), .B0(\key_mem[0][84] ), .B1(n5761), 
        .Y(n1781) );
  AO22X1 U3414 ( .A0(n4014), .A1(n1510), .B0(\key_mem[14][85] ), .B1(n4024), 
        .Y(n3572) );
  AO22X1 U3415 ( .A0(n4070), .A1(n1510), .B0(\key_mem[12][85] ), .B1(n4079), 
        .Y(n3316) );
  AO22X1 U3416 ( .A0(n4126), .A1(n1510), .B0(\key_mem[10][85] ), .B1(n4134), 
        .Y(n3060) );
  AO22X1 U3417 ( .A0(n4182), .A1(n1510), .B0(\key_mem[8][85] ), .B1(n4190), 
        .Y(n2804) );
  AO22X1 U3418 ( .A0(n4239), .A1(n1510), .B0(\key_mem[6][85] ), .B1(n4252), 
        .Y(n2548) );
  AO22X1 U3419 ( .A0(n4294), .A1(n1510), .B0(\key_mem[4][85] ), .B1(n4300), 
        .Y(n2292) );
  AO22X1 U3420 ( .A0(n4350), .A1(n1510), .B0(\key_mem[2][85] ), .B1(n4363), 
        .Y(n2036) );
  AO22X1 U3421 ( .A0(n3951), .A1(n1510), .B0(\key_mem[0][85] ), .B1(n5761), 
        .Y(n1780) );
  AO22X1 U3422 ( .A0(n4014), .A1(n1512), .B0(\key_mem[14][87] ), .B1(n4022), 
        .Y(n3570) );
  AO22X1 U3423 ( .A0(n4070), .A1(n1512), .B0(\key_mem[12][87] ), .B1(n4078), 
        .Y(n3314) );
  AO22X1 U3424 ( .A0(n4126), .A1(n1512), .B0(\key_mem[10][87] ), .B1(n4133), 
        .Y(n3058) );
  AO22X1 U3425 ( .A0(n4182), .A1(n1512), .B0(\key_mem[8][87] ), .B1(n4189), 
        .Y(n2802) );
  AO22X1 U3426 ( .A0(n4239), .A1(n1512), .B0(\key_mem[6][87] ), .B1(n4251), 
        .Y(n2546) );
  AO22X1 U3427 ( .A0(n4294), .A1(n1512), .B0(\key_mem[4][87] ), .B1(n4299), 
        .Y(n2290) );
  AO22X1 U3428 ( .A0(n4350), .A1(n1512), .B0(\key_mem[2][87] ), .B1(n4362), 
        .Y(n2034) );
  AO22X1 U3429 ( .A0(n3951), .A1(n1512), .B0(\key_mem[0][87] ), .B1(n5761), 
        .Y(n1778) );
  AO22X1 U3430 ( .A0(n4015), .A1(n1522), .B0(\key_mem[14][97] ), .B1(n4022), 
        .Y(n3560) );
  AO22X1 U3431 ( .A0(n4071), .A1(n1522), .B0(\key_mem[12][97] ), .B1(n4078), 
        .Y(n3304) );
  AO22X1 U3432 ( .A0(n4127), .A1(n1522), .B0(\key_mem[10][97] ), .B1(n4140), 
        .Y(n3048) );
  AO22X1 U3433 ( .A0(n4183), .A1(n1522), .B0(\key_mem[8][97] ), .B1(n4196), 
        .Y(n2792) );
  AO22X1 U3434 ( .A0(n4240), .A1(n1522), .B0(\key_mem[6][97] ), .B1(n4252), 
        .Y(n2536) );
  AO22X1 U3435 ( .A0(n4295), .A1(n1522), .B0(\key_mem[4][97] ), .B1(n4302), 
        .Y(n2280) );
  AO22X1 U3436 ( .A0(n4351), .A1(n1522), .B0(\key_mem[2][97] ), .B1(n4362), 
        .Y(n2024) );
  AO22X1 U3437 ( .A0(n3950), .A1(n1522), .B0(\key_mem[0][97] ), .B1(n3932), 
        .Y(n1768) );
  AO22X1 U3438 ( .A0(n4015), .A1(n1523), .B0(\key_mem[14][98] ), .B1(n4021), 
        .Y(n3559) );
  AO22X1 U3439 ( .A0(n4071), .A1(n1523), .B0(\key_mem[12][98] ), .B1(n4077), 
        .Y(n3303) );
  AO22X1 U3440 ( .A0(n4127), .A1(n1523), .B0(\key_mem[10][98] ), .B1(n4142), 
        .Y(n3047) );
  AO22X1 U3441 ( .A0(n4183), .A1(n1523), .B0(\key_mem[8][98] ), .B1(n4198), 
        .Y(n2791) );
  AO22X1 U3442 ( .A0(n4240), .A1(n1523), .B0(\key_mem[6][98] ), .B1(n4251), 
        .Y(n2535) );
  AO22X1 U3443 ( .A0(n4295), .A1(n1523), .B0(\key_mem[4][98] ), .B1(n4301), 
        .Y(n2279) );
  AO22X1 U3444 ( .A0(n4351), .A1(n1523), .B0(\key_mem[2][98] ), .B1(n4359), 
        .Y(n2023) );
  AO22X1 U3445 ( .A0(n3950), .A1(n1523), .B0(\key_mem[0][98] ), .B1(n3932), 
        .Y(n1767) );
  AO22X1 U3446 ( .A0(n4015), .A1(n1524), .B0(\key_mem[14][99] ), .B1(n4020), 
        .Y(n3558) );
  AO22X1 U3447 ( .A0(n4071), .A1(n1524), .B0(\key_mem[12][99] ), .B1(n4076), 
        .Y(n3302) );
  AO22X1 U3448 ( .A0(n4127), .A1(n1524), .B0(\key_mem[10][99] ), .B1(n4141), 
        .Y(n3046) );
  AO22X1 U3449 ( .A0(n4183), .A1(n1524), .B0(\key_mem[8][99] ), .B1(n4197), 
        .Y(n2790) );
  AO22X1 U3450 ( .A0(n4240), .A1(n1524), .B0(\key_mem[6][99] ), .B1(n4248), 
        .Y(n2534) );
  AO22X1 U3451 ( .A0(n4295), .A1(n1524), .B0(\key_mem[4][99] ), .B1(n4300), 
        .Y(n2278) );
  AO22X1 U3452 ( .A0(n4351), .A1(n1524), .B0(\key_mem[2][99] ), .B1(n4358), 
        .Y(n2022) );
  AO22X1 U3453 ( .A0(n3950), .A1(n1524), .B0(\key_mem[0][99] ), .B1(n1717), 
        .Y(n1766) );
  AO22X1 U3454 ( .A0(n4016), .A1(n1525), .B0(\key_mem[14][100] ), .B1(n4019), 
        .Y(n3557) );
  AO22X1 U3455 ( .A0(n4072), .A1(n1525), .B0(\key_mem[12][100] ), .B1(n4075), 
        .Y(n3301) );
  AO22X1 U3456 ( .A0(n4128), .A1(n1525), .B0(\key_mem[10][100] ), .B1(n4140), 
        .Y(n3045) );
  AO22X1 U3457 ( .A0(n4184), .A1(n1525), .B0(\key_mem[8][100] ), .B1(n4196), 
        .Y(n2789) );
  AO22X1 U3458 ( .A0(n4241), .A1(n1525), .B0(\key_mem[6][100] ), .B1(n4247), 
        .Y(n2533) );
  AO22X1 U3459 ( .A0(n4296), .A1(n1525), .B0(\key_mem[4][100] ), .B1(n4299), 
        .Y(n2277) );
  AO22X1 U3460 ( .A0(n4352), .A1(n1525), .B0(\key_mem[2][100] ), .B1(n4357), 
        .Y(n2021) );
  AO22X1 U3461 ( .A0(n3950), .A1(n1525), .B0(\key_mem[0][100] ), .B1(n1717), 
        .Y(n1765) );
  AO22X1 U3462 ( .A0(n4016), .A1(n1526), .B0(\key_mem[14][101] ), .B1(n4026), 
        .Y(n3556) );
  AO22X1 U3463 ( .A0(n4072), .A1(n1526), .B0(\key_mem[12][101] ), .B1(n4087), 
        .Y(n3300) );
  AO22X1 U3464 ( .A0(n4128), .A1(n1526), .B0(\key_mem[10][101] ), .B1(n4142), 
        .Y(n3044) );
  AO22X1 U3465 ( .A0(n4184), .A1(n1526), .B0(\key_mem[8][101] ), .B1(n4198), 
        .Y(n2788) );
  AO22X1 U3466 ( .A0(n4241), .A1(n1526), .B0(\key_mem[6][101] ), .B1(n4246), 
        .Y(n2532) );
  AO22X1 U3467 ( .A0(n4296), .A1(n1526), .B0(\key_mem[4][101] ), .B1(n4304), 
        .Y(n2276) );
  AO22X1 U3468 ( .A0(n4352), .A1(n1526), .B0(\key_mem[2][101] ), .B1(n4356), 
        .Y(n2020) );
  AO22X1 U3469 ( .A0(n3950), .A1(n1526), .B0(\key_mem[0][101] ), .B1(n1717), 
        .Y(n1764) );
  AO22X1 U3470 ( .A0(n4016), .A1(n1528), .B0(\key_mem[14][103] ), .B1(n4029), 
        .Y(n3554) );
  AO22X1 U3471 ( .A0(n4072), .A1(n1528), .B0(\key_mem[12][103] ), .B1(n4084), 
        .Y(n3298) );
  AO22X1 U3472 ( .A0(n4128), .A1(n1528), .B0(\key_mem[10][103] ), .B1(n4136), 
        .Y(n3042) );
  AO22X1 U3473 ( .A0(n4184), .A1(n1528), .B0(\key_mem[8][103] ), .B1(n4192), 
        .Y(n2786) );
  AO22X1 U3474 ( .A0(n4241), .A1(n1528), .B0(\key_mem[6][103] ), .B1(n4247), 
        .Y(n2530) );
  AO22X1 U3475 ( .A0(n4296), .A1(n1528), .B0(\key_mem[4][103] ), .B1(n4308), 
        .Y(n2274) );
  AO22X1 U3476 ( .A0(n4352), .A1(n1528), .B0(\key_mem[2][103] ), .B1(n4355), 
        .Y(n2018) );
  AO22X1 U3477 ( .A0(n3949), .A1(n1528), .B0(\key_mem[0][103] ), .B1(n1717), 
        .Y(n1762) );
  AO22X1 U3478 ( .A0(n4016), .A1(n1530), .B0(\key_mem[14][105] ), .B1(n740), 
        .Y(n3552) );
  AO22X1 U3479 ( .A0(n4072), .A1(n1530), .B0(\key_mem[12][105] ), .B1(n4084), 
        .Y(n3296) );
  AO22X1 U3480 ( .A0(n4128), .A1(n1530), .B0(\key_mem[10][105] ), .B1(n4135), 
        .Y(n3040) );
  AO22X1 U3481 ( .A0(n4184), .A1(n1530), .B0(\key_mem[8][105] ), .B1(n4191), 
        .Y(n2784) );
  AO22X1 U3482 ( .A0(n4241), .A1(n1530), .B0(\key_mem[6][105] ), .B1(n4253), 
        .Y(n2528) );
  AO22X1 U3483 ( .A0(n4296), .A1(n1530), .B0(\key_mem[4][105] ), .B1(n4300), 
        .Y(n2272) );
  AO22X1 U3484 ( .A0(n4352), .A1(n1530), .B0(\key_mem[2][105] ), .B1(n4359), 
        .Y(n2016) );
  AO22X1 U3485 ( .A0(n3949), .A1(n1530), .B0(\key_mem[0][105] ), .B1(n1717), 
        .Y(n1760) );
  AO22X1 U3486 ( .A0(n4016), .A1(n1531), .B0(\key_mem[14][106] ), .B1(n4026), 
        .Y(n3551) );
  AO22X1 U3487 ( .A0(n4072), .A1(n1531), .B0(\key_mem[12][106] ), .B1(n4084), 
        .Y(n3295) );
  AO22X1 U3488 ( .A0(n4128), .A1(n1531), .B0(\key_mem[10][106] ), .B1(n4134), 
        .Y(n3039) );
  AO22X1 U3489 ( .A0(n4184), .A1(n1531), .B0(\key_mem[8][106] ), .B1(n4190), 
        .Y(n2783) );
  AO22X1 U3490 ( .A0(n4241), .A1(n1531), .B0(\key_mem[6][106] ), .B1(n4254), 
        .Y(n2527) );
  AO22X1 U3491 ( .A0(n4296), .A1(n1531), .B0(\key_mem[4][106] ), .B1(n4304), 
        .Y(n2271) );
  AO22X1 U3492 ( .A0(n4352), .A1(n1531), .B0(\key_mem[2][106] ), .B1(n4365), 
        .Y(n2015) );
  AO22X1 U3493 ( .A0(n3949), .A1(n1531), .B0(\key_mem[0][106] ), .B1(n1717), 
        .Y(n1759) );
  AO22X1 U3494 ( .A0(n4016), .A1(n1533), .B0(\key_mem[14][108] ), .B1(n4025), 
        .Y(n3549) );
  AO22X1 U3495 ( .A0(n4072), .A1(n1533), .B0(\key_mem[12][108] ), .B1(n4084), 
        .Y(n3293) );
  AO22X1 U3496 ( .A0(n4128), .A1(n1533), .B0(\key_mem[10][108] ), .B1(n4133), 
        .Y(n3037) );
  AO22X1 U3497 ( .A0(n4184), .A1(n1533), .B0(\key_mem[8][108] ), .B1(n4189), 
        .Y(n2781) );
  AO22X1 U3498 ( .A0(n4241), .A1(n1533), .B0(\key_mem[6][108] ), .B1(n4250), 
        .Y(n2525) );
  AO22X1 U3499 ( .A0(n4296), .A1(n1533), .B0(\key_mem[4][108] ), .B1(n4303), 
        .Y(n2269) );
  AO22X1 U3500 ( .A0(n4352), .A1(n1533), .B0(\key_mem[2][108] ), .B1(n4364), 
        .Y(n2013) );
  AO22X1 U3501 ( .A0(n3949), .A1(n1533), .B0(\key_mem[0][108] ), .B1(n1717), 
        .Y(n1757) );
  AO22X1 U3502 ( .A0(n4016), .A1(n1534), .B0(\key_mem[14][109] ), .B1(n4023), 
        .Y(n3548) );
  AO22X1 U3503 ( .A0(n4072), .A1(n1534), .B0(\key_mem[12][109] ), .B1(n4084), 
        .Y(n3292) );
  AO22X1 U3504 ( .A0(n4128), .A1(n1534), .B0(\key_mem[10][109] ), .B1(n4139), 
        .Y(n3036) );
  AO22X1 U3505 ( .A0(n4184), .A1(n1534), .B0(\key_mem[8][109] ), .B1(n4195), 
        .Y(n2780) );
  AO22X1 U3506 ( .A0(n4241), .A1(n1534), .B0(\key_mem[6][109] ), .B1(n4254), 
        .Y(n2524) );
  AO22X1 U3507 ( .A0(n4296), .A1(n1534), .B0(\key_mem[4][109] ), .B1(n4302), 
        .Y(n2268) );
  AO22X1 U3508 ( .A0(n4352), .A1(n1534), .B0(\key_mem[2][109] ), .B1(n4363), 
        .Y(n2012) );
  AO22X1 U3509 ( .A0(n3949), .A1(n1534), .B0(\key_mem[0][109] ), .B1(n3933), 
        .Y(n1756) );
  AO22X1 U3510 ( .A0(n4017), .A1(n1536), .B0(\key_mem[14][111] ), .B1(n4024), 
        .Y(n3546) );
  AO22X1 U3511 ( .A0(n4073), .A1(n1536), .B0(\key_mem[12][111] ), .B1(n4084), 
        .Y(n3290) );
  AO22X1 U3512 ( .A0(n4129), .A1(n1536), .B0(\key_mem[10][111] ), .B1(n4138), 
        .Y(n3034) );
  AO22X1 U3513 ( .A0(n4185), .A1(n1536), .B0(\key_mem[8][111] ), .B1(n4194), 
        .Y(n2778) );
  AO22X1 U3514 ( .A0(n4242), .A1(n1536), .B0(\key_mem[6][111] ), .B1(n4247), 
        .Y(n2522) );
  AO22X1 U3515 ( .A0(n4297), .A1(n1536), .B0(\key_mem[4][111] ), .B1(n4301), 
        .Y(n2266) );
  AO22X1 U3516 ( .A0(n4353), .A1(n1536), .B0(\key_mem[2][111] ), .B1(n4362), 
        .Y(n2010) );
  AO22X1 U3517 ( .A0(n3949), .A1(n1536), .B0(\key_mem[0][111] ), .B1(n3933), 
        .Y(n1754) );
  AO22X1 U3518 ( .A0(n4017), .A1(n1537), .B0(\key_mem[14][112] ), .B1(n4022), 
        .Y(n3545) );
  AO22X1 U3519 ( .A0(n4073), .A1(n1537), .B0(\key_mem[12][112] ), .B1(n4084), 
        .Y(n3289) );
  AO22X1 U3520 ( .A0(n4129), .A1(n1537), .B0(\key_mem[10][112] ), .B1(n4137), 
        .Y(n3033) );
  AO22X1 U3521 ( .A0(n4185), .A1(n1537), .B0(\key_mem[8][112] ), .B1(n4193), 
        .Y(n2777) );
  AO22X1 U3522 ( .A0(n4242), .A1(n1537), .B0(\key_mem[6][112] ), .B1(n4254), 
        .Y(n2521) );
  AO22X1 U3523 ( .A0(n4297), .A1(n1537), .B0(\key_mem[4][112] ), .B1(n4300), 
        .Y(n2265) );
  AO22X1 U3524 ( .A0(n4353), .A1(n1537), .B0(\key_mem[2][112] ), .B1(n4361), 
        .Y(n2009) );
  AO22X1 U3525 ( .A0(n3949), .A1(n1537), .B0(\key_mem[0][112] ), .B1(n3933), 
        .Y(n1753) );
  AO22X1 U3526 ( .A0(n4017), .A1(n1538), .B0(\key_mem[14][113] ), .B1(n4023), 
        .Y(n3544) );
  AO22X1 U3527 ( .A0(n4073), .A1(n1538), .B0(\key_mem[12][113] ), .B1(n4085), 
        .Y(n3288) );
  AO22X1 U3528 ( .A0(n4129), .A1(n1538), .B0(\key_mem[10][113] ), .B1(n4139), 
        .Y(n3032) );
  AO22X1 U3529 ( .A0(n4185), .A1(n1538), .B0(\key_mem[8][113] ), .B1(n4195), 
        .Y(n2776) );
  AO22X1 U3530 ( .A0(n4242), .A1(n1538), .B0(\key_mem[6][113] ), .B1(n4246), 
        .Y(n2520) );
  AO22X1 U3531 ( .A0(n4297), .A1(n1538), .B0(\key_mem[4][113] ), .B1(n4309), 
        .Y(n2264) );
  AO22X1 U3532 ( .A0(n4353), .A1(n1538), .B0(\key_mem[2][113] ), .B1(n4362), 
        .Y(n2008) );
  AO22X1 U3533 ( .A0(n3948), .A1(n1538), .B0(\key_mem[0][113] ), .B1(n3933), 
        .Y(n1752) );
  AO22X1 U3534 ( .A0(n4017), .A1(n1539), .B0(\key_mem[14][114] ), .B1(n4024), 
        .Y(n3543) );
  AO22X1 U3535 ( .A0(n4073), .A1(n1539), .B0(\key_mem[12][114] ), .B1(n4085), 
        .Y(n3287) );
  AO22X1 U3536 ( .A0(n4129), .A1(n1539), .B0(\key_mem[10][114] ), .B1(n4138), 
        .Y(n3031) );
  AO22X1 U3537 ( .A0(n4185), .A1(n1539), .B0(\key_mem[8][114] ), .B1(n4194), 
        .Y(n2775) );
  AO22X1 U3538 ( .A0(n4242), .A1(n1539), .B0(\key_mem[6][114] ), .B1(n4245), 
        .Y(n2519) );
  AO22X1 U3539 ( .A0(n4297), .A1(n1539), .B0(\key_mem[4][114] ), .B1(n4308), 
        .Y(n2263) );
  AO22X1 U3540 ( .A0(n4353), .A1(n1539), .B0(\key_mem[2][114] ), .B1(n4361), 
        .Y(n2007) );
  AO22X1 U3541 ( .A0(n3948), .A1(n1539), .B0(\key_mem[0][114] ), .B1(n3933), 
        .Y(n1751) );
  AO22X1 U3542 ( .A0(n4017), .A1(n1541), .B0(\key_mem[14][116] ), .B1(n4022), 
        .Y(n3541) );
  AO22X1 U3543 ( .A0(n4073), .A1(n1541), .B0(\key_mem[12][116] ), .B1(n4085), 
        .Y(n3285) );
  AO22X1 U3544 ( .A0(n4129), .A1(n1541), .B0(\key_mem[10][116] ), .B1(n4137), 
        .Y(n3029) );
  AO22X1 U3545 ( .A0(n4185), .A1(n1541), .B0(\key_mem[8][116] ), .B1(n4193), 
        .Y(n2773) );
  AO22X1 U3546 ( .A0(n4242), .A1(n1541), .B0(\key_mem[6][116] ), .B1(n4254), 
        .Y(n2517) );
  AO22X1 U3547 ( .A0(n4297), .A1(n1541), .B0(\key_mem[4][116] ), .B1(n4309), 
        .Y(n2261) );
  AO22X1 U3548 ( .A0(n4353), .A1(n1541), .B0(\key_mem[2][116] ), .B1(n4360), 
        .Y(n2005) );
  AO22X1 U3549 ( .A0(n3948), .A1(n1541), .B0(\key_mem[0][116] ), .B1(n3933), 
        .Y(n1749) );
  AO22X1 U3550 ( .A0(n4017), .A1(n1542), .B0(\key_mem[14][117] ), .B1(n4021), 
        .Y(n3540) );
  AO22X1 U3551 ( .A0(n4073), .A1(n1542), .B0(\key_mem[12][117] ), .B1(n4085), 
        .Y(n3284) );
  AO22X1 U3552 ( .A0(n4129), .A1(n1542), .B0(\key_mem[10][117] ), .B1(n4140), 
        .Y(n3028) );
  AO22X1 U3553 ( .A0(n4185), .A1(n1542), .B0(\key_mem[8][117] ), .B1(n4196), 
        .Y(n2772) );
  AO22X1 U3554 ( .A0(n4242), .A1(n1542), .B0(\key_mem[6][117] ), .B1(n4245), 
        .Y(n2516) );
  AO22X1 U3555 ( .A0(n4297), .A1(n1542), .B0(\key_mem[4][117] ), .B1(n4308), 
        .Y(n2260) );
  AO22X1 U3556 ( .A0(n4353), .A1(n1542), .B0(\key_mem[2][117] ), .B1(n4359), 
        .Y(n2004) );
  AO22X1 U3557 ( .A0(n3948), .A1(n1542), .B0(\key_mem[0][117] ), .B1(n3933), 
        .Y(n1748) );
  AO22X1 U3558 ( .A0(n4017), .A1(n1543), .B0(\key_mem[14][118] ), .B1(n4020), 
        .Y(n3539) );
  AO22X1 U3559 ( .A0(n4073), .A1(n1543), .B0(\key_mem[12][118] ), .B1(n4085), 
        .Y(n3283) );
  AO22X1 U3560 ( .A0(n4129), .A1(n1543), .B0(\key_mem[10][118] ), .B1(n4131), 
        .Y(n3027) );
  AO22X1 U3561 ( .A0(n4185), .A1(n1543), .B0(\key_mem[8][118] ), .B1(n4187), 
        .Y(n2771) );
  AO22X1 U3562 ( .A0(n4242), .A1(n1543), .B0(\key_mem[6][118] ), .B1(n4253), 
        .Y(n2515) );
  AO22X1 U3563 ( .A0(n4297), .A1(n1543), .B0(\key_mem[4][118] ), .B1(n4309), 
        .Y(n2259) );
  AO22X1 U3564 ( .A0(n4353), .A1(n1543), .B0(\key_mem[2][118] ), .B1(n4358), 
        .Y(n2003) );
  AO22X1 U3565 ( .A0(n3948), .A1(n1543), .B0(\key_mem[0][118] ), .B1(n3933), 
        .Y(n1747) );
  AO22X1 U3566 ( .A0(n4017), .A1(n1544), .B0(\key_mem[14][119] ), .B1(n4019), 
        .Y(n3538) );
  AO22X1 U3567 ( .A0(n4073), .A1(n1544), .B0(\key_mem[12][119] ), .B1(n4085), 
        .Y(n3282) );
  AO22X1 U3568 ( .A0(n4129), .A1(n1544), .B0(\key_mem[10][119] ), .B1(n4132), 
        .Y(n3026) );
  AO22X1 U3569 ( .A0(n4185), .A1(n1544), .B0(\key_mem[8][119] ), .B1(n4188), 
        .Y(n2770) );
  AO22X1 U3570 ( .A0(n4242), .A1(n1544), .B0(\key_mem[6][119] ), .B1(n4254), 
        .Y(n2514) );
  AO22X1 U3571 ( .A0(n4297), .A1(n1544), .B0(\key_mem[4][119] ), .B1(n4308), 
        .Y(n2258) );
  AO22X1 U3572 ( .A0(n4353), .A1(n1544), .B0(\key_mem[2][119] ), .B1(n4363), 
        .Y(n2002) );
  AO22X1 U3573 ( .A0(n3948), .A1(n1544), .B0(\key_mem[0][119] ), .B1(n3934), 
        .Y(n1746) );
  AO22X1 U3574 ( .A0(n3968), .A1(n1474), .B0(\key_mem[1][49] ), .B1(n5762), 
        .Y(n1944) );
  AO22X1 U3575 ( .A0(n4038), .A1(n1474), .B0(\key_mem[13][49] ), .B1(n4047), 
        .Y(n3480) );
  AO22X1 U3576 ( .A0(n4094), .A1(n671), .B0(\key_mem[11][49] ), .B1(n4104), 
        .Y(n3224) );
  AO22X1 U3577 ( .A0(n4150), .A1(n671), .B0(\key_mem[9][49] ), .B1(n4160), .Y(
        n2968) );
  AO22X1 U3578 ( .A0(n4202), .A1(n671), .B0(\key_mem[7][49] ), .B1(n4217), .Y(
        n2712) );
  AO22X1 U3579 ( .A0(n4262), .A1(n671), .B0(\key_mem[5][49] ), .B1(n4271), .Y(
        n2456) );
  AO22X1 U3580 ( .A0(n4318), .A1(n671), .B0(\key_mem[3][49] ), .B1(n4340), .Y(
        n2200) );
  AO22X1 U3581 ( .A0(n4010), .A1(n1474), .B0(\key_mem[14][49] ), .B1(n4019), 
        .Y(n3608) );
  AO22X1 U3582 ( .A0(n4066), .A1(n1474), .B0(\key_mem[12][49] ), .B1(n4080), 
        .Y(n3352) );
  AO22X1 U3583 ( .A0(n4122), .A1(n1474), .B0(\key_mem[10][49] ), .B1(n4141), 
        .Y(n3096) );
  AO22X1 U3584 ( .A0(n4178), .A1(n1474), .B0(\key_mem[8][49] ), .B1(n4197), 
        .Y(n2840) );
  AO22X1 U3585 ( .A0(n4235), .A1(n1474), .B0(\key_mem[6][49] ), .B1(n4257), 
        .Y(n2584) );
  AO22X1 U3586 ( .A0(n4290), .A1(n1474), .B0(\key_mem[4][49] ), .B1(n4310), 
        .Y(n2328) );
  AO22X1 U3587 ( .A0(n4346), .A1(n1474), .B0(\key_mem[2][49] ), .B1(n4360), 
        .Y(n2072) );
  AO22X1 U3588 ( .A0(n3955), .A1(n1474), .B0(\key_mem[0][49] ), .B1(n3928), 
        .Y(n1816) );
  AO22X1 U3589 ( .A0(n3966), .A1(n1445), .B0(\key_mem[1][20] ), .B1(n3991), 
        .Y(n1973) );
  AO22X1 U3590 ( .A0(n3969), .A1(n1479), .B0(\key_mem[1][54] ), .B1(n5762), 
        .Y(n1939) );
  AO22X1 U3591 ( .A0(n4036), .A1(n1445), .B0(\key_mem[13][20] ), .B1(n4056), 
        .Y(n3509) );
  AO22X1 U3592 ( .A0(n4092), .A1(n700), .B0(\key_mem[11][20] ), .B1(n4110), 
        .Y(n3253) );
  AO22X1 U3593 ( .A0(n4148), .A1(n700), .B0(\key_mem[9][20] ), .B1(n4163), .Y(
        n2997) );
  AO22X1 U3594 ( .A0(n4205), .A1(n700), .B0(\key_mem[7][20] ), .B1(n4221), .Y(
        n2741) );
  AO22X1 U3595 ( .A0(n4260), .A1(n700), .B0(\key_mem[5][20] ), .B1(n4275), .Y(
        n2485) );
  AO22X1 U3596 ( .A0(n4316), .A1(n700), .B0(\key_mem[3][20] ), .B1(n4340), .Y(
        n2229) );
  AO22X1 U3597 ( .A0(n4039), .A1(n1479), .B0(\key_mem[13][54] ), .B1(n4058), 
        .Y(n3475) );
  AO22X1 U3598 ( .A0(n4095), .A1(n666), .B0(\key_mem[11][54] ), .B1(n4116), 
        .Y(n3219) );
  AO22X1 U3599 ( .A0(n4151), .A1(n666), .B0(\key_mem[9][54] ), .B1(n4168), .Y(
        n2963) );
  AO22X1 U3600 ( .A0(n4207), .A1(n666), .B0(\key_mem[7][54] ), .B1(n4219), .Y(
        n2707) );
  AO22X1 U3601 ( .A0(n4263), .A1(n666), .B0(\key_mem[5][54] ), .B1(n4282), .Y(
        n2451) );
  AO22X1 U3602 ( .A0(n4319), .A1(n666), .B0(\key_mem[3][54] ), .B1(n4329), .Y(
        n2195) );
  AO22X1 U3603 ( .A0(n3965), .A1(n1437), .B0(\key_mem[1][12] ), .B1(n3981), 
        .Y(n1981) );
  AO22X1 U3604 ( .A0(n3959), .A1(n1434), .B0(\key_mem[0][9] ), .B1(n1719), .Y(
        n1856) );
  AO22X1 U3605 ( .A0(n4035), .A1(n1437), .B0(\key_mem[13][12] ), .B1(n4052), 
        .Y(n3517) );
  AO22X1 U3606 ( .A0(n4091), .A1(n708), .B0(\key_mem[11][12] ), .B1(n4114), 
        .Y(n3261) );
  AO22X1 U3607 ( .A0(n4147), .A1(n708), .B0(\key_mem[9][12] ), .B1(n4170), .Y(
        n3005) );
  AO22X1 U3608 ( .A0(n4204), .A1(n708), .B0(\key_mem[7][12] ), .B1(n4220), .Y(
        n2749) );
  AO22X1 U3609 ( .A0(n4259), .A1(n708), .B0(\key_mem[5][12] ), .B1(n4282), .Y(
        n2493) );
  AO22X1 U3610 ( .A0(n4315), .A1(n708), .B0(\key_mem[3][12] ), .B1(n4330), .Y(
        n2237) );
  AO22X1 U3611 ( .A0(n3959), .A1(n1437), .B0(\key_mem[0][12] ), .B1(n1720), 
        .Y(n1853) );
  AO22X1 U3612 ( .A0(n3958), .A1(n1441), .B0(\key_mem[0][16] ), .B1(n1720), 
        .Y(n1849) );
  AO22X1 U3613 ( .A0(n3958), .A1(n1442), .B0(\key_mem[0][17] ), .B1(n1720), 
        .Y(n1848) );
  AO22X1 U3614 ( .A0(n3958), .A1(n1445), .B0(\key_mem[0][20] ), .B1(n1720), 
        .Y(n1845) );
  AO22X1 U3615 ( .A0(n3972), .A1(n1505), .B0(\key_mem[1][80] ), .B1(n3978), 
        .Y(n1913) );
  AO22X1 U3616 ( .A0(n3972), .A1(n1511), .B0(\key_mem[1][86] ), .B1(n3977), 
        .Y(n1907) );
  AO22X1 U3617 ( .A0(n4042), .A1(n1505), .B0(\key_mem[13][80] ), .B1(n4048), 
        .Y(n3449) );
  AO22X1 U3618 ( .A0(n4098), .A1(n640), .B0(\key_mem[11][80] ), .B1(n4114), 
        .Y(n3193) );
  AO22X1 U3619 ( .A0(n4154), .A1(n640), .B0(\key_mem[9][80] ), .B1(n4165), .Y(
        n2937) );
  AO22X1 U3620 ( .A0(n4210), .A1(n640), .B0(\key_mem[7][80] ), .B1(n4216), .Y(
        n2681) );
  AO22X1 U3621 ( .A0(n4266), .A1(n640), .B0(\key_mem[5][80] ), .B1(n4278), .Y(
        n2425) );
  AO22X1 U3622 ( .A0(n4322), .A1(n640), .B0(\key_mem[3][80] ), .B1(n4332), .Y(
        n2169) );
  AO22X1 U3623 ( .A0(n4042), .A1(n1511), .B0(\key_mem[13][86] ), .B1(n4061), 
        .Y(n3443) );
  AO22X1 U3624 ( .A0(n4098), .A1(n1511), .B0(\key_mem[11][86] ), .B1(n4103), 
        .Y(n3187) );
  AO22X1 U3625 ( .A0(n4154), .A1(n1511), .B0(\key_mem[9][86] ), .B1(n4160), 
        .Y(n2931) );
  AO22X1 U3626 ( .A0(n4210), .A1(n1511), .B0(\key_mem[7][86] ), .B1(n4228), 
        .Y(n2675) );
  AO22X1 U3627 ( .A0(n4266), .A1(n1511), .B0(\key_mem[5][86] ), .B1(n4279), 
        .Y(n2419) );
  AO22X1 U3628 ( .A0(n4322), .A1(n1511), .B0(\key_mem[3][86] ), .B1(n4332), 
        .Y(n2163) );
  AO22X1 U3629 ( .A0(n3964), .A1(n1434), .B0(\key_mem[1][9] ), .B1(n3983), .Y(
        n1984) );
  AO22X1 U3630 ( .A0(n3965), .A1(n1441), .B0(\key_mem[1][16] ), .B1(n3979), 
        .Y(n1977) );
  AO22X1 U3631 ( .A0(n3965), .A1(n1442), .B0(\key_mem[1][17] ), .B1(n3986), 
        .Y(n1976) );
  AO22X1 U3632 ( .A0(n3968), .A1(n1466), .B0(\key_mem[1][41] ), .B1(n3982), 
        .Y(n1952) );
  AO22X1 U3633 ( .A0(n3968), .A1(n1469), .B0(\key_mem[1][44] ), .B1(n3985), 
        .Y(n1949) );
  AO22X1 U3634 ( .A0(n3969), .A1(n1477), .B0(\key_mem[1][52] ), .B1(n5762), 
        .Y(n1941) );
  AO22X1 U3635 ( .A0(n3971), .A1(n1498), .B0(\key_mem[1][73] ), .B1(n3983), 
        .Y(n1920) );
  AO22X1 U3636 ( .A0(n3971), .A1(n1501), .B0(\key_mem[1][76] ), .B1(n3982), 
        .Y(n1917) );
  AO22X1 U3637 ( .A0(n4007), .A1(n1441), .B0(\key_mem[14][16] ), .B1(n4032), 
        .Y(n3641) );
  AO22X1 U3638 ( .A0(n4035), .A1(n1441), .B0(\key_mem[13][16] ), .B1(n4055), 
        .Y(n3513) );
  AO22X1 U3639 ( .A0(n4063), .A1(n1441), .B0(\key_mem[12][16] ), .B1(n4075), 
        .Y(n3385) );
  AO22X1 U3640 ( .A0(n4091), .A1(n1441), .B0(\key_mem[11][16] ), .B1(n4113), 
        .Y(n3257) );
  AO22X1 U3641 ( .A0(n4119), .A1(n704), .B0(\key_mem[10][16] ), .B1(n4138), 
        .Y(n3129) );
  AO22X1 U3642 ( .A0(n4147), .A1(n1441), .B0(\key_mem[9][16] ), .B1(n4160), 
        .Y(n3001) );
  AO22X1 U3643 ( .A0(n4175), .A1(n704), .B0(\key_mem[8][16] ), .B1(n4194), .Y(
        n2873) );
  AO22X1 U3644 ( .A0(n4204), .A1(n1441), .B0(\key_mem[7][16] ), .B1(n4221), 
        .Y(n2745) );
  AO22X1 U3645 ( .A0(n4232), .A1(n704), .B0(\key_mem[6][16] ), .B1(n4248), .Y(
        n2617) );
  AO22X1 U3646 ( .A0(n4259), .A1(n1441), .B0(\key_mem[5][16] ), .B1(n4279), 
        .Y(n2489) );
  AO22X1 U3647 ( .A0(n4287), .A1(n704), .B0(\key_mem[4][16] ), .B1(n4313), .Y(
        n2361) );
  AO22X1 U3648 ( .A0(n4315), .A1(n1441), .B0(\key_mem[3][16] ), .B1(n4337), 
        .Y(n2233) );
  AO22X1 U3649 ( .A0(n4343), .A1(n704), .B0(\key_mem[2][16] ), .B1(n4362), .Y(
        n2105) );
  AO22X1 U3650 ( .A0(n4007), .A1(n1442), .B0(\key_mem[14][17] ), .B1(n4023), 
        .Y(n3640) );
  AO22X1 U3651 ( .A0(n4063), .A1(n1442), .B0(\key_mem[12][17] ), .B1(n4079), 
        .Y(n3384) );
  AO22X1 U3652 ( .A0(n4119), .A1(n703), .B0(\key_mem[10][17] ), .B1(n4131), 
        .Y(n3128) );
  AO22X1 U3653 ( .A0(n4175), .A1(n703), .B0(\key_mem[8][17] ), .B1(n4187), .Y(
        n2872) );
  AO22X1 U3654 ( .A0(n4232), .A1(n703), .B0(\key_mem[6][17] ), .B1(n4255), .Y(
        n2616) );
  AO22X1 U3655 ( .A0(n4287), .A1(n703), .B0(\key_mem[4][17] ), .B1(n4304), .Y(
        n2360) );
  AO22X1 U3656 ( .A0(n4343), .A1(n703), .B0(\key_mem[2][17] ), .B1(n4365), .Y(
        n2104) );
  AO22X1 U3657 ( .A0(n4008), .A1(n1445), .B0(\key_mem[14][20] ), .B1(n4022), 
        .Y(n3637) );
  AO22X1 U3658 ( .A0(n4064), .A1(n1445), .B0(\key_mem[12][20] ), .B1(n4088), 
        .Y(n3381) );
  AO22X1 U3659 ( .A0(n4120), .A1(n1445), .B0(\key_mem[10][20] ), .B1(n736), 
        .Y(n3125) );
  AO22X1 U3660 ( .A0(n4176), .A1(n1445), .B0(\key_mem[8][20] ), .B1(n733), .Y(
        n2869) );
  AO22X1 U3661 ( .A0(n4233), .A1(n1445), .B0(\key_mem[6][20] ), .B1(n4252), 
        .Y(n2613) );
  AO22X1 U3662 ( .A0(n4288), .A1(n1445), .B0(\key_mem[4][20] ), .B1(n4313), 
        .Y(n2357) );
  AO22X1 U3663 ( .A0(n4344), .A1(n1445), .B0(\key_mem[2][20] ), .B1(n4359), 
        .Y(n2101) );
  AO22X1 U3664 ( .A0(n4010), .A1(n1466), .B0(\key_mem[14][41] ), .B1(n4028), 
        .Y(n3616) );
  AO22X1 U3665 ( .A0(n4038), .A1(n1466), .B0(\key_mem[13][41] ), .B1(n4061), 
        .Y(n3488) );
  AO22X1 U3666 ( .A0(n4066), .A1(n1466), .B0(\key_mem[12][41] ), .B1(n4087), 
        .Y(n3360) );
  AO22X1 U3667 ( .A0(n4094), .A1(n679), .B0(\key_mem[11][41] ), .B1(n4103), 
        .Y(n3232) );
  AO22X1 U3668 ( .A0(n4122), .A1(n1466), .B0(\key_mem[10][41] ), .B1(n4138), 
        .Y(n3104) );
  AO22X1 U3669 ( .A0(n4150), .A1(n679), .B0(\key_mem[9][41] ), .B1(n4163), .Y(
        n2976) );
  AO22X1 U3670 ( .A0(n4178), .A1(n1466), .B0(\key_mem[8][41] ), .B1(n4194), 
        .Y(n2848) );
  AO22X1 U3671 ( .A0(n4202), .A1(n679), .B0(\key_mem[7][41] ), .B1(n4223), .Y(
        n2720) );
  AO22X1 U3672 ( .A0(n4235), .A1(n1466), .B0(\key_mem[6][41] ), .B1(n4244), 
        .Y(n2592) );
  AO22X1 U3673 ( .A0(n4262), .A1(n679), .B0(\key_mem[5][41] ), .B1(n4274), .Y(
        n2464) );
  AO22X1 U3674 ( .A0(n4290), .A1(n1466), .B0(\key_mem[4][41] ), .B1(n4301), 
        .Y(n2336) );
  AO22X1 U3675 ( .A0(n4318), .A1(n679), .B0(\key_mem[3][41] ), .B1(n4335), .Y(
        n2208) );
  AO22X1 U3676 ( .A0(n4346), .A1(n1466), .B0(\key_mem[2][41] ), .B1(n4369), 
        .Y(n2080) );
  AO22X1 U3677 ( .A0(n3956), .A1(n1466), .B0(\key_mem[0][41] ), .B1(n3928), 
        .Y(n1824) );
  AO22X1 U3678 ( .A0(n4010), .A1(n1469), .B0(\key_mem[14][44] ), .B1(n4030), 
        .Y(n3613) );
  AO22X1 U3679 ( .A0(n4038), .A1(n1469), .B0(\key_mem[13][44] ), .B1(n4054), 
        .Y(n3485) );
  AO22X1 U3680 ( .A0(n4066), .A1(n1469), .B0(\key_mem[12][44] ), .B1(n4079), 
        .Y(n3357) );
  AO22X1 U3681 ( .A0(n4094), .A1(n676), .B0(\key_mem[11][44] ), .B1(n4110), 
        .Y(n3229) );
  AO22X1 U3682 ( .A0(n4122), .A1(n1469), .B0(\key_mem[10][44] ), .B1(n4136), 
        .Y(n3101) );
  AO22X1 U3683 ( .A0(n4150), .A1(n676), .B0(\key_mem[9][44] ), .B1(n4167), .Y(
        n2973) );
  AO22X1 U3684 ( .A0(n4178), .A1(n1469), .B0(\key_mem[8][44] ), .B1(n4190), 
        .Y(n2845) );
  AO22X1 U3685 ( .A0(n4202), .A1(n676), .B0(\key_mem[7][44] ), .B1(n4220), .Y(
        n2717) );
  AO22X1 U3686 ( .A0(n4235), .A1(n1469), .B0(\key_mem[6][44] ), .B1(n4257), 
        .Y(n2589) );
  AO22X1 U3687 ( .A0(n4262), .A1(n676), .B0(\key_mem[5][44] ), .B1(n4278), .Y(
        n2461) );
  AO22X1 U3688 ( .A0(n4290), .A1(n1469), .B0(\key_mem[4][44] ), .B1(n4299), 
        .Y(n2333) );
  AO22X1 U3689 ( .A0(n4318), .A1(n676), .B0(\key_mem[3][44] ), .B1(n4338), .Y(
        n2205) );
  AO22X1 U3690 ( .A0(n4346), .A1(n1469), .B0(\key_mem[2][44] ), .B1(n4355), 
        .Y(n2077) );
  AO22X1 U3691 ( .A0(n3955), .A1(n1469), .B0(\key_mem[0][44] ), .B1(n3928), 
        .Y(n1821) );
  AO22X1 U3692 ( .A0(n4011), .A1(n1477), .B0(\key_mem[14][52] ), .B1(n4028), 
        .Y(n3605) );
  AO22X1 U3693 ( .A0(n4039), .A1(n1477), .B0(\key_mem[13][52] ), .B1(n4048), 
        .Y(n3477) );
  AO22X1 U3694 ( .A0(n4067), .A1(n1477), .B0(\key_mem[12][52] ), .B1(n4078), 
        .Y(n3349) );
  AO22X1 U3695 ( .A0(n4095), .A1(n668), .B0(\key_mem[11][52] ), .B1(n4111), 
        .Y(n3221) );
  AO22X1 U3696 ( .A0(n4123), .A1(n1477), .B0(\key_mem[10][52] ), .B1(n4136), 
        .Y(n3093) );
  AO22X1 U3697 ( .A0(n4151), .A1(n668), .B0(\key_mem[9][52] ), .B1(n4162), .Y(
        n2965) );
  AO22X1 U3698 ( .A0(n4179), .A1(n1477), .B0(\key_mem[8][52] ), .B1(n4192), 
        .Y(n2837) );
  AO22X1 U3699 ( .A0(n4207), .A1(n668), .B0(\key_mem[7][52] ), .B1(n4219), .Y(
        n2709) );
  AO22X1 U3700 ( .A0(n4236), .A1(n1477), .B0(\key_mem[6][52] ), .B1(n4257), 
        .Y(n2581) );
  AO22X1 U3701 ( .A0(n4263), .A1(n668), .B0(\key_mem[5][52] ), .B1(n4278), .Y(
        n2453) );
  AO22X1 U3702 ( .A0(n4291), .A1(n1477), .B0(\key_mem[4][52] ), .B1(n4311), 
        .Y(n2325) );
  AO22X1 U3703 ( .A0(n4319), .A1(n668), .B0(\key_mem[3][52] ), .B1(n4333), .Y(
        n2197) );
  AO22X1 U3704 ( .A0(n4347), .A1(n1477), .B0(\key_mem[2][52] ), .B1(n4367), 
        .Y(n2069) );
  AO22X1 U3705 ( .A0(n3955), .A1(n1477), .B0(\key_mem[0][52] ), .B1(n3929), 
        .Y(n1813) );
  AO22X1 U3706 ( .A0(n4011), .A1(n1479), .B0(\key_mem[14][54] ), .B1(n4024), 
        .Y(n3603) );
  AO22X1 U3707 ( .A0(n4067), .A1(n1479), .B0(\key_mem[12][54] ), .B1(n4076), 
        .Y(n3347) );
  AO22X1 U3708 ( .A0(n4123), .A1(n1479), .B0(\key_mem[10][54] ), .B1(n4133), 
        .Y(n3091) );
  AO22X1 U3709 ( .A0(n4179), .A1(n1479), .B0(\key_mem[8][54] ), .B1(n4189), 
        .Y(n2835) );
  AO22X1 U3710 ( .A0(n4236), .A1(n1479), .B0(\key_mem[6][54] ), .B1(n4247), 
        .Y(n2579) );
  AO22X1 U3711 ( .A0(n4291), .A1(n1479), .B0(\key_mem[4][54] ), .B1(n727), .Y(
        n2323) );
  AO22X1 U3712 ( .A0(n4347), .A1(n1479), .B0(\key_mem[2][54] ), .B1(n4355), 
        .Y(n2067) );
  AO22X1 U3713 ( .A0(n3954), .A1(n1479), .B0(\key_mem[0][54] ), .B1(n3929), 
        .Y(n1811) );
  AO22X1 U3714 ( .A0(n4013), .A1(n1498), .B0(\key_mem[14][73] ), .B1(n4019), 
        .Y(n3584) );
  AO22X1 U3715 ( .A0(n4041), .A1(n1498), .B0(\key_mem[13][73] ), .B1(n4056), 
        .Y(n3456) );
  AO22X1 U3716 ( .A0(n4069), .A1(n1498), .B0(\key_mem[12][73] ), .B1(n4083), 
        .Y(n3328) );
  AO22X1 U3717 ( .A0(n4097), .A1(n647), .B0(\key_mem[11][73] ), .B1(n4104), 
        .Y(n3200) );
  AO22X1 U3718 ( .A0(n4125), .A1(n1498), .B0(\key_mem[10][73] ), .B1(n4135), 
        .Y(n3072) );
  AO22X1 U3719 ( .A0(n4153), .A1(n647), .B0(\key_mem[9][73] ), .B1(n4166), .Y(
        n2944) );
  AO22X1 U3720 ( .A0(n4181), .A1(n1498), .B0(\key_mem[8][73] ), .B1(n4192), 
        .Y(n2816) );
  AO22X1 U3721 ( .A0(n4209), .A1(n647), .B0(\key_mem[7][73] ), .B1(n4215), .Y(
        n2688) );
  AO22X1 U3722 ( .A0(n4238), .A1(n1498), .B0(\key_mem[6][73] ), .B1(n4247), 
        .Y(n2560) );
  AO22X1 U3723 ( .A0(n4265), .A1(n647), .B0(\key_mem[5][73] ), .B1(n4272), .Y(
        n2432) );
  AO22X1 U3724 ( .A0(n4293), .A1(n1498), .B0(\key_mem[4][73] ), .B1(n4300), 
        .Y(n2304) );
  AO22X1 U3725 ( .A0(n4321), .A1(n647), .B0(\key_mem[3][73] ), .B1(n4331), .Y(
        n2176) );
  AO22X1 U3726 ( .A0(n4349), .A1(n1498), .B0(\key_mem[2][73] ), .B1(n4366), 
        .Y(n2048) );
  AO22X1 U3727 ( .A0(n3952), .A1(n1498), .B0(\key_mem[0][73] ), .B1(n3931), 
        .Y(n1792) );
  AO22X1 U3728 ( .A0(n4013), .A1(n1501), .B0(\key_mem[14][76] ), .B1(n4022), 
        .Y(n3581) );
  AO22X1 U3729 ( .A0(n4041), .A1(n1501), .B0(\key_mem[13][76] ), .B1(n4055), 
        .Y(n3453) );
  AO22X1 U3730 ( .A0(n4069), .A1(n1501), .B0(\key_mem[12][76] ), .B1(n4082), 
        .Y(n3325) );
  AO22X1 U3731 ( .A0(n4097), .A1(n644), .B0(\key_mem[11][76] ), .B1(n4103), 
        .Y(n3197) );
  AO22X1 U3732 ( .A0(n4125), .A1(n1501), .B0(\key_mem[10][76] ), .B1(n4134), 
        .Y(n3069) );
  AO22X1 U3733 ( .A0(n4153), .A1(n644), .B0(\key_mem[9][76] ), .B1(n4159), .Y(
        n2941) );
  AO22X1 U3734 ( .A0(n4181), .A1(n1501), .B0(\key_mem[8][76] ), .B1(n4191), 
        .Y(n2813) );
  AO22X1 U3735 ( .A0(n4209), .A1(n644), .B0(\key_mem[7][76] ), .B1(n4228), .Y(
        n2685) );
  AO22X1 U3736 ( .A0(n4238), .A1(n1501), .B0(\key_mem[6][76] ), .B1(n4246), 
        .Y(n2557) );
  AO22X1 U3737 ( .A0(n4265), .A1(n644), .B0(\key_mem[5][76] ), .B1(n4271), .Y(
        n2429) );
  AO22X1 U3738 ( .A0(n4293), .A1(n1501), .B0(\key_mem[4][76] ), .B1(n4299), 
        .Y(n2301) );
  AO22X1 U3739 ( .A0(n4321), .A1(n644), .B0(\key_mem[3][76] ), .B1(n4329), .Y(
        n2173) );
  AO22X1 U3740 ( .A0(n4349), .A1(n1501), .B0(\key_mem[2][76] ), .B1(n4366), 
        .Y(n2045) );
  AO22X1 U3741 ( .A0(n3952), .A1(n1501), .B0(\key_mem[0][76] ), .B1(n3931), 
        .Y(n1789) );
  AO22X1 U3742 ( .A0(n4014), .A1(n1505), .B0(\key_mem[14][80] ), .B1(n4026), 
        .Y(n3577) );
  AO22X1 U3743 ( .A0(n4070), .A1(n1505), .B0(\key_mem[12][80] ), .B1(n4081), 
        .Y(n3321) );
  AO22X1 U3744 ( .A0(n4126), .A1(n1505), .B0(\key_mem[10][80] ), .B1(n4133), 
        .Y(n3065) );
  AO22X1 U3745 ( .A0(n4182), .A1(n1505), .B0(\key_mem[8][80] ), .B1(n4189), 
        .Y(n2809) );
  AO22X1 U3746 ( .A0(n4239), .A1(n1505), .B0(\key_mem[6][80] ), .B1(n4247), 
        .Y(n2553) );
  AO22X1 U3747 ( .A0(n4294), .A1(n1505), .B0(\key_mem[4][80] ), .B1(n4304), 
        .Y(n2297) );
  AO22X1 U3748 ( .A0(n4350), .A1(n1505), .B0(\key_mem[2][80] ), .B1(n4366), 
        .Y(n2041) );
  AO22X1 U3749 ( .A0(n3952), .A1(n1505), .B0(\key_mem[0][80] ), .B1(n5761), 
        .Y(n1785) );
  AO22X1 U3750 ( .A0(n4014), .A1(n1511), .B0(\key_mem[14][86] ), .B1(n4021), 
        .Y(n3571) );
  AO22X1 U3751 ( .A0(n4070), .A1(n1511), .B0(\key_mem[12][86] ), .B1(n4077), 
        .Y(n3315) );
  AO22X1 U3752 ( .A0(n4126), .A1(n1511), .B0(\key_mem[10][86] ), .B1(n4131), 
        .Y(n3059) );
  AO22X1 U3753 ( .A0(n4182), .A1(n634), .B0(\key_mem[8][86] ), .B1(n4187), .Y(
        n2803) );
  AO22X1 U3754 ( .A0(n4239), .A1(n634), .B0(\key_mem[6][86] ), .B1(n4250), .Y(
        n2547) );
  AO22X1 U3755 ( .A0(n4294), .A1(n634), .B0(\key_mem[4][86] ), .B1(n4304), .Y(
        n2291) );
  AO22X1 U3756 ( .A0(n4350), .A1(n634), .B0(\key_mem[2][86] ), .B1(n4361), .Y(
        n2035) );
  AO22X1 U3757 ( .A0(n3951), .A1(n634), .B0(\key_mem[0][86] ), .B1(n5761), .Y(
        n1779) );
  AO22X1 U3758 ( .A0(n4007), .A1(n1437), .B0(\key_mem[14][12] ), .B1(n4029), 
        .Y(n3645) );
  AO22X1 U3759 ( .A0(n4063), .A1(n1437), .B0(\key_mem[12][12] ), .B1(n738), 
        .Y(n3389) );
  AO22X1 U3760 ( .A0(n4119), .A1(n1437), .B0(\key_mem[10][12] ), .B1(n4142), 
        .Y(n3133) );
  AO22X1 U3761 ( .A0(n4175), .A1(n1437), .B0(\key_mem[8][12] ), .B1(n4198), 
        .Y(n2877) );
  AO22X1 U3762 ( .A0(n4232), .A1(n1437), .B0(\key_mem[6][12] ), .B1(n4253), 
        .Y(n2621) );
  AO22X1 U3763 ( .A0(n4287), .A1(n1437), .B0(\key_mem[4][12] ), .B1(n4303), 
        .Y(n2365) );
  AO22X1 U3764 ( .A0(n4343), .A1(n1437), .B0(\key_mem[2][12] ), .B1(n4360), 
        .Y(n2109) );
  AO22X1 U3765 ( .A0(n4006), .A1(n1434), .B0(\key_mem[14][9] ), .B1(n4026), 
        .Y(n3648) );
  AO22X1 U3766 ( .A0(n4034), .A1(n1434), .B0(\key_mem[13][9] ), .B1(n4055), 
        .Y(n3520) );
  AO22X1 U3767 ( .A0(n4062), .A1(n1434), .B0(\key_mem[12][9] ), .B1(n4083), 
        .Y(n3392) );
  AO22X1 U3768 ( .A0(n4090), .A1(n711), .B0(\key_mem[11][9] ), .B1(n4111), .Y(
        n3264) );
  AO22X1 U3769 ( .A0(n4118), .A1(n1434), .B0(\key_mem[10][9] ), .B1(n4139), 
        .Y(n3136) );
  AO22X1 U3770 ( .A0(n4146), .A1(n711), .B0(\key_mem[9][9] ), .B1(n4167), .Y(
        n3008) );
  AO22X1 U3771 ( .A0(n4174), .A1(n1434), .B0(\key_mem[8][9] ), .B1(n4195), .Y(
        n2880) );
  AO22X1 U3772 ( .A0(n4203), .A1(n711), .B0(\key_mem[7][9] ), .B1(n4217), .Y(
        n2752) );
  AO22X1 U3773 ( .A0(n4231), .A1(n1434), .B0(\key_mem[6][9] ), .B1(n4252), .Y(
        n2624) );
  AO22X1 U3774 ( .A0(n4258), .A1(n711), .B0(\key_mem[5][9] ), .B1(n4279), .Y(
        n2496) );
  AO22X1 U3775 ( .A0(n4286), .A1(n1434), .B0(\key_mem[4][9] ), .B1(n4307), .Y(
        n2368) );
  AO22X1 U3776 ( .A0(n4314), .A1(n711), .B0(\key_mem[3][9] ), .B1(n4335), .Y(
        n2240) );
  AO22X1 U3777 ( .A0(n4342), .A1(n1434), .B0(\key_mem[2][9] ), .B1(n4363), .Y(
        n2112) );
  XNOR2X1 U3778 ( .A(n5266), .B(prev_key1_reg[84]), .Y(n32) );
  AO22X1 U3779 ( .A0(prev_key1_reg[127]), .A1(n1616), .B0(n1602), .B1(n5636), 
        .Y(n5637) );
  INVX1 U3780 ( .A(n741), .Y(n5636) );
  XNOR2X1 U3781 ( .A(n5014), .B(sboxw[12]), .Y(n33) );
  AO22X1 U3782 ( .A0(sboxw[16]), .A1(n1610), .B0(n1597), .B1(n5148), .Y(n5149)
         );
  AO22X1 U3783 ( .A0(sboxw[17]), .A1(n1611), .B0(n1598), .B1(n5181), .Y(n5182)
         );
  AO22X1 U3784 ( .A0(sboxw[22]), .A1(n1613), .B0(n1600), .B1(n5345), .Y(n5346)
         );
  AO22X1 U3785 ( .A0(prev_key1_reg[48]), .A1(n1610), .B0(n1597), .B1(n5136), 
        .Y(n5137) );
  AO22X1 U3786 ( .A0(prev_key1_reg[49]), .A1(n1611), .B0(n1598), .B1(n5169), 
        .Y(n5170) );
  AO22X1 U3787 ( .A0(prev_key1_reg[80]), .A1(n1610), .B0(n1597), .B1(n5128), 
        .Y(n5129) );
  AO22X1 U3788 ( .A0(prev_key1_reg[81]), .A1(n1610), .B0(n1597), .B1(n5161), 
        .Y(n5162) );
  AO22X1 U3789 ( .A0(prev_key1_reg[86]), .A1(n1612), .B0(n1599), .B1(n5326), 
        .Y(n5327) );
  XNOR2X1 U3790 ( .A(n4743), .B(prev_key1_reg[68]), .Y(n34) );
  XNOR2X1 U3791 ( .A(n4616), .B(prev_key1_reg[64]), .Y(n35) );
  XNOR2X1 U3792 ( .A(n4754), .B(sboxw[4]), .Y(n36) );
  AO22X1 U3793 ( .A0(sboxw[18]), .A1(n1611), .B0(n1598), .B1(n5214), .Y(n5215)
         );
  AO22X1 U3794 ( .A0(sboxw[19]), .A1(n1611), .B0(n1598), .B1(n5247), .Y(n5248)
         );
  AO22X1 U3795 ( .A0(sboxw[21]), .A1(n1612), .B0(n1599), .B1(n5313), .Y(n5314)
         );
  AO22X1 U3796 ( .A0(sboxw[23]), .A1(n1613), .B0(n1600), .B1(n5378), .Y(n5379)
         );
  AO22X1 U3797 ( .A0(prev_key1_reg[50]), .A1(n1611), .B0(n1598), .B1(n5202), 
        .Y(n5203) );
  AO22X1 U3798 ( .A0(prev_key1_reg[51]), .A1(n1611), .B0(n1598), .B1(n5235), 
        .Y(n5236) );
  AO22X1 U3799 ( .A0(prev_key1_reg[53]), .A1(n1612), .B0(n1599), .B1(n5301), 
        .Y(n5302) );
  AO22X1 U3800 ( .A0(prev_key1_reg[55]), .A1(n1613), .B0(n1600), .B1(n5366), 
        .Y(n5367) );
  AO22X1 U3801 ( .A0(prev_key1_reg[82]), .A1(n1611), .B0(n1598), .B1(n5194), 
        .Y(n5195) );
  AO22X1 U3802 ( .A0(prev_key1_reg[83]), .A1(n1611), .B0(n1598), .B1(n5227), 
        .Y(n5228) );
  AO22X1 U3803 ( .A0(prev_key1_reg[85]), .A1(n1612), .B0(n1599), .B1(n5293), 
        .Y(n5294) );
  AO22X1 U3804 ( .A0(prev_key1_reg[87]), .A1(n1613), .B0(n1600), .B1(n5358), 
        .Y(n5359) );
  XNOR2X1 U3805 ( .A(n4679), .B(prev_key1_reg[66]), .Y(n37) );
  XNOR2X1 U3806 ( .A(n4711), .B(prev_key1_reg[67]), .Y(n38) );
  XNOR2X1 U3807 ( .A(n4775), .B(prev_key1_reg[69]), .Y(n39) );
  XNOR2X1 U3808 ( .A(n4806), .B(prev_key1_reg[70]), .Y(n40) );
  XNOR2X1 U3809 ( .A(n4838), .B(prev_key1_reg[71]), .Y(n41) );
  XNOR2X1 U3810 ( .A(n4937), .B(prev_key1_reg[74]), .Y(n42) );
  XNOR2X1 U3811 ( .A(n4970), .B(prev_key1_reg[75]), .Y(n43) );
  XNOR2X1 U3812 ( .A(n5036), .B(prev_key1_reg[77]), .Y(n44) );
  XNOR2X1 U3813 ( .A(n5101), .B(prev_key1_reg[79]), .Y(n45) );
  XNOR2X1 U3814 ( .A(n5200), .B(prev_key1_reg[82]), .Y(n46) );
  XNOR2X1 U3815 ( .A(n5299), .B(prev_key1_reg[85]), .Y(n47) );
  XNOR2X1 U3816 ( .A(n5364), .B(prev_key1_reg[87]), .Y(n48) );
  XNOR2X1 U3817 ( .A(n4626), .B(sboxw[0]), .Y(n49) );
  XNOR2X1 U3818 ( .A(n4690), .B(sboxw[2]), .Y(n50) );
  XNOR2X1 U3819 ( .A(n4722), .B(sboxw[3]), .Y(n51) );
  XNOR2X1 U3820 ( .A(n4786), .B(sboxw[5]), .Y(n52) );
  XNOR2X1 U3821 ( .A(n4817), .B(sboxw[6]), .Y(n53) );
  XNOR2X1 U3822 ( .A(n4849), .B(sboxw[7]), .Y(n54) );
  XNOR2X1 U3823 ( .A(n4948), .B(sboxw[10]), .Y(n55) );
  XNOR2X1 U3824 ( .A(n4981), .B(sboxw[11]), .Y(n56) );
  XNOR2X1 U3825 ( .A(n5047), .B(sboxw[13]), .Y(n57) );
  XNOR2X1 U3826 ( .A(n5211), .B(sboxw[18]), .Y(n58) );
  XNOR2X1 U3827 ( .A(n5447), .B(prev_key1_reg[121]), .Y(n59) );
  XNOR2X1 U3828 ( .A(n5555), .B(prev_key1_reg[124]), .Y(n60) );
  XNOR2X1 U3829 ( .A(n5591), .B(prev_key1_reg[125]), .Y(n61) );
  XNOR2X1 U3830 ( .A(n5627), .B(prev_key1_reg[126]), .Y(n62) );
  XNOR2X1 U3831 ( .A(n5519), .B(prev_key1_reg[123]), .Y(n63) );
  XNOR2X1 U3832 ( .A(n5483), .B(prev_key1_reg[122]), .Y(n64) );
  XNOR2X1 U3833 ( .A(n5411), .B(prev_key1_reg[120]), .Y(n65) );
  XNOR2X1 U3834 ( .A(n5134), .B(prev_key1_reg[80]), .Y(n66) );
  XNOR2X1 U3835 ( .A(n5167), .B(prev_key1_reg[81]), .Y(n67) );
  XNOR2X1 U3836 ( .A(n5332), .B(prev_key1_reg[86]), .Y(n68) );
  XNOR2X1 U3837 ( .A(n5003), .B(prev_key1_reg[76]), .Y(n69) );
  XNOR2X1 U3838 ( .A(n4915), .B(sboxw[9]), .Y(n70) );
  XNOR2X1 U3839 ( .A(n5145), .B(sboxw[16]), .Y(n71) );
  XNOR2X1 U3840 ( .A(n5178), .B(sboxw[17]), .Y(n72) );
  XNOR2X1 U3841 ( .A(n5277), .B(sboxw[20]), .Y(n73) );
  XNOR2X1 U3842 ( .A(n5342), .B(sboxw[22]), .Y(n74) );
  AO22X1 U3843 ( .A0(sboxw[31]), .A1(n1616), .B0(n1602), .B1(n5667), .Y(n5670)
         );
  INVX1 U3844 ( .A(n1129), .Y(n5667) );
  AO22X1 U3845 ( .A0(prev_key1_reg[63]), .A1(n1616), .B0(n1604), .B1(n5653), 
        .Y(n5654) );
  INVX1 U3846 ( .A(n1001), .Y(n5653) );
  AO22X1 U3847 ( .A0(prev_key1_reg[95]), .A1(n1616), .B0(n1604), .B1(n5644), 
        .Y(n5645) );
  INVX1 U3848 ( .A(n873), .Y(n5644) );
  AO22X1 U3849 ( .A0(n672), .A1(n4094), .B0(\key_mem[11][48] ), .B1(n4114), 
        .Y(n3225) );
  AO22X1 U3850 ( .A0(n4315), .A1(n1442), .B0(\key_mem[3][17] ), .B1(n4334), 
        .Y(n2232) );
  AO22X1 U3851 ( .A0(n4259), .A1(n1442), .B0(\key_mem[5][17] ), .B1(n729), .Y(
        n2488) );
  AO22X1 U3852 ( .A0(n4204), .A1(n1442), .B0(\key_mem[7][17] ), .B1(n4221), 
        .Y(n2744) );
  AO22X1 U3853 ( .A0(n4147), .A1(n1442), .B0(\key_mem[9][17] ), .B1(n735), .Y(
        n3000) );
  AO22X1 U3854 ( .A0(n4091), .A1(n1442), .B0(\key_mem[11][17] ), .B1(n4111), 
        .Y(n3256) );
  AO22X1 U3855 ( .A0(n4035), .A1(n1442), .B0(\key_mem[13][17] ), .B1(n4054), 
        .Y(n3512) );
  AO22X1 U3856 ( .A0(n4038), .A1(n1473), .B0(\key_mem[13][48] ), .B1(n4061), 
        .Y(n3481) );
  AO22X1 U3857 ( .A0(n4150), .A1(n1473), .B0(\key_mem[9][48] ), .B1(n4165), 
        .Y(n2969) );
  AO22X1 U3858 ( .A0(n4202), .A1(n672), .B0(\key_mem[7][48] ), .B1(n4218), .Y(
        n2713) );
  AO22X1 U3859 ( .A0(n4262), .A1(n672), .B0(\key_mem[5][48] ), .B1(n4272), .Y(
        n2457) );
  AO22X1 U3860 ( .A0(n4318), .A1(n672), .B0(\key_mem[3][48] ), .B1(n4327), .Y(
        n2201) );
  AO22X1 U3861 ( .A0(n3968), .A1(n672), .B0(\key_mem[1][48] ), .B1(n5762), .Y(
        n1945) );
  AO22X1 U3862 ( .A0(n3955), .A1(n1473), .B0(\key_mem[0][48] ), .B1(n3928), 
        .Y(n1817) );
  AO22X1 U3863 ( .A0(n4346), .A1(n1473), .B0(\key_mem[2][48] ), .B1(n4368), 
        .Y(n2073) );
  AO22X1 U3864 ( .A0(n4290), .A1(n1473), .B0(\key_mem[4][48] ), .B1(n4312), 
        .Y(n2329) );
  AO22X1 U3865 ( .A0(n4235), .A1(n1473), .B0(\key_mem[6][48] ), .B1(n4257), 
        .Y(n2585) );
  AO22X1 U3866 ( .A0(n4178), .A1(n1473), .B0(\key_mem[8][48] ), .B1(n4192), 
        .Y(n2841) );
  AO22X1 U3867 ( .A0(n4122), .A1(n1473), .B0(\key_mem[10][48] ), .B1(n4135), 
        .Y(n3097) );
  AO22X1 U3868 ( .A0(n4066), .A1(n1473), .B0(\key_mem[12][48] ), .B1(n4077), 
        .Y(n3353) );
  AO22X1 U3869 ( .A0(n4010), .A1(n1473), .B0(\key_mem[14][48] ), .B1(n4032), 
        .Y(n3609) );
  OAI221XL U3870 ( .A0(n1667), .A1(n4896), .B0(n4895), .B1(n1657), .C0(n4894), 
        .Y(n3807) );
  INVX1 U3871 ( .A(key[105]), .Y(n4896) );
  AOI221XL U3872 ( .A0(n1646), .A1(n835), .B0(n1631), .B1(key[233]), .C0(n4893), .Y(n4894) );
  AO22X1 U3873 ( .A0(prev_key1_reg[105]), .A1(n1620), .B0(n1607), .B1(n4892), 
        .Y(n4893) );
  OAI221XL U3874 ( .A0(n1672), .A1(n5454), .B0(n5453), .B1(n1655), .C0(n5452), 
        .Y(n3887) );
  INVX1 U3875 ( .A(key[25]), .Y(n5454) );
  AOI221XL U3876 ( .A0(n1649), .A1(n24), .B0(n1630), .B1(key[153]), .C0(n5451), 
        .Y(n5452) );
  AO22X1 U3877 ( .A0(sboxw[25]), .A1(n1614), .B0(n1601), .B1(n5450), .Y(n5451)
         );
  OAI221XL U3878 ( .A0(n1672), .A1(n5441), .B0(n5440), .B1(n1655), .C0(n5439), 
        .Y(n3855) );
  INVX1 U3879 ( .A(key[57]), .Y(n5441) );
  AOI221XL U3880 ( .A0(n1646), .A1(n17), .B0(n1630), .B1(key[185]), .C0(n5438), 
        .Y(n5439) );
  AO22X1 U3881 ( .A0(prev_key1_reg[57]), .A1(n1614), .B0(n1601), .B1(n5437), 
        .Y(n5438) );
  OAI221XL U3882 ( .A0(n1672), .A1(n5431), .B0(n5430), .B1(n1655), .C0(n5429), 
        .Y(n3823) );
  INVX1 U3883 ( .A(key[89]), .Y(n5431) );
  AOI221XL U3884 ( .A0(n1648), .A1(n899), .B0(n1630), .B1(key[217]), .C0(n5428), .Y(n5429) );
  AO22X1 U3885 ( .A0(prev_key1_reg[89]), .A1(n1614), .B0(n1601), .B1(n5427), 
        .Y(n5428) );
  OAI221XL U3886 ( .A0(n1664), .A1(n5562), .B0(n5561), .B1(n1653), .C0(n5560), 
        .Y(n3884) );
  INVX1 U3887 ( .A(key[28]), .Y(n5562) );
  AOI221XL U3888 ( .A0(n1648), .A1(n25), .B0(n1635), .B1(key[156]), .C0(n5559), 
        .Y(n5560) );
  AO22X1 U3889 ( .A0(sboxw[28]), .A1(n1615), .B0(n1602), .B1(n5558), .Y(n5559)
         );
  OAI221XL U3890 ( .A0(n1677), .A1(n5549), .B0(n5548), .B1(n1653), .C0(n5547), 
        .Y(n3852) );
  INVX1 U3891 ( .A(key[60]), .Y(n5549) );
  AOI221XL U3892 ( .A0(n1647), .A1(n18), .B0(n1633), .B1(key[188]), .C0(n5546), 
        .Y(n5547) );
  AO22X1 U3893 ( .A0(prev_key1_reg[60]), .A1(n1615), .B0(n1607), .B1(n5545), 
        .Y(n5546) );
  OAI221XL U3894 ( .A0(n1674), .A1(n5539), .B0(n5538), .B1(n1653), .C0(n5537), 
        .Y(n3820) );
  INVX1 U3895 ( .A(key[92]), .Y(n5539) );
  AOI221XL U3896 ( .A0(n1648), .A1(n887), .B0(n1633), .B1(key[220]), .C0(n5536), .Y(n5537) );
  AO22X1 U3897 ( .A0(prev_key1_reg[92]), .A1(n1615), .B0(n1602), .B1(n5535), 
        .Y(n5536) );
  OAI221XL U3898 ( .A0(n1675), .A1(n5598), .B0(n5597), .B1(n1655), .C0(n5596), 
        .Y(n3883) );
  INVX1 U3899 ( .A(key[29]), .Y(n5598) );
  AOI221XL U3900 ( .A0(n1636), .A1(n26), .B0(n1631), .B1(key[157]), .C0(n5595), 
        .Y(n5596) );
  AO22X1 U3901 ( .A0(sboxw[29]), .A1(n1615), .B0(n1603), .B1(n5594), .Y(n5595)
         );
  OAI221XL U3902 ( .A0(n1676), .A1(n5585), .B0(n5584), .B1(n1654), .C0(n5583), 
        .Y(n3851) );
  INVX1 U3903 ( .A(key[61]), .Y(n5585) );
  AOI221XL U3904 ( .A0(n1636), .A1(n19), .B0(n5671), .B1(key[189]), .C0(n5582), 
        .Y(n5583) );
  AO22X1 U3905 ( .A0(prev_key1_reg[61]), .A1(n1615), .B0(n1605), .B1(n5581), 
        .Y(n5582) );
  OAI221XL U3906 ( .A0(n1673), .A1(n5575), .B0(n5574), .B1(n1653), .C0(n5573), 
        .Y(n3819) );
  INVX1 U3907 ( .A(key[93]), .Y(n5575) );
  AOI221XL U3908 ( .A0(n1648), .A1(n883), .B0(n1634), .B1(key[221]), .C0(n5572), .Y(n5573) );
  AO22X1 U3909 ( .A0(prev_key1_reg[93]), .A1(n1615), .B0(n1602), .B1(n5571), 
        .Y(n5572) );
  OAI221XL U3910 ( .A0(n1676), .A1(n5634), .B0(n5633), .B1(n1654), .C0(n5632), 
        .Y(n3882) );
  INVX1 U3911 ( .A(key[30]), .Y(n5634) );
  AOI221XL U3912 ( .A0(n1636), .A1(n27), .B0(n5671), .B1(key[158]), .C0(n5631), 
        .Y(n5632) );
  AO22X1 U3913 ( .A0(sboxw[30]), .A1(n1616), .B0(n1605), .B1(n5630), .Y(n5631)
         );
  OAI221XL U3914 ( .A0(n1664), .A1(n5621), .B0(n5620), .B1(n1653), .C0(n5619), 
        .Y(n3850) );
  INVX1 U3915 ( .A(key[62]), .Y(n5621) );
  AOI221XL U3916 ( .A0(n1636), .A1(n20), .B0(n1635), .B1(key[190]), .C0(n5618), 
        .Y(n5619) );
  AO22X1 U3917 ( .A0(prev_key1_reg[62]), .A1(n1616), .B0(n1607), .B1(n5617), 
        .Y(n5618) );
  OAI221XL U3918 ( .A0(n1674), .A1(n5611), .B0(n5610), .B1(n1654), .C0(n5609), 
        .Y(n3818) );
  INVX1 U3919 ( .A(key[94]), .Y(n5611) );
  AOI221XL U3920 ( .A0(n1636), .A1(n879), .B0(n1632), .B1(key[222]), .C0(n5608), .Y(n5609) );
  AO22X1 U3921 ( .A0(prev_key1_reg[94]), .A1(n1616), .B0(n1602), .B1(n5607), 
        .Y(n5608) );
  OAI221XL U3922 ( .A0(n1677), .A1(n5526), .B0(n5525), .B1(n1655), .C0(n5524), 
        .Y(n3885) );
  INVX1 U3923 ( .A(key[27]), .Y(n5526) );
  AOI221XL U3924 ( .A0(n1645), .A1(n28), .B0(n5671), .B1(key[155]), .C0(n5523), 
        .Y(n5524) );
  AO22X1 U3925 ( .A0(sboxw[27]), .A1(n1615), .B0(n1604), .B1(n5522), .Y(n5523)
         );
  OAI221XL U3926 ( .A0(n1675), .A1(n5513), .B0(n5512), .B1(n1653), .C0(n5511), 
        .Y(n3853) );
  INVX1 U3927 ( .A(key[59]), .Y(n5513) );
  AOI221XL U3928 ( .A0(n1649), .A1(n21), .B0(n5671), .B1(key[187]), .C0(n5510), 
        .Y(n5511) );
  AO22X1 U3929 ( .A0(prev_key1_reg[59]), .A1(n1615), .B0(n1607), .B1(n5509), 
        .Y(n5510) );
  OAI221XL U3930 ( .A0(n1672), .A1(n5503), .B0(n5502), .B1(n1654), .C0(n5501), 
        .Y(n3821) );
  INVX1 U3931 ( .A(key[91]), .Y(n5503) );
  AOI221XL U3932 ( .A0(n1648), .A1(n891), .B0(n1630), .B1(key[219]), .C0(n5500), .Y(n5501) );
  AO22X1 U3933 ( .A0(prev_key1_reg[91]), .A1(n1614), .B0(n1601), .B1(n5499), 
        .Y(n5500) );
  OAI221XL U3934 ( .A0(n1672), .A1(n5490), .B0(n5489), .B1(n1654), .C0(n5488), 
        .Y(n3886) );
  INVX1 U3935 ( .A(key[26]), .Y(n5490) );
  AOI221XL U3936 ( .A0(n1647), .A1(n29), .B0(n1630), .B1(key[154]), .C0(n5487), 
        .Y(n5488) );
  AO22X1 U3937 ( .A0(sboxw[26]), .A1(n1614), .B0(n1601), .B1(n5486), .Y(n5487)
         );
  OAI221XL U3938 ( .A0(n1672), .A1(n5477), .B0(n5476), .B1(n1655), .C0(n5475), 
        .Y(n3854) );
  INVX1 U3939 ( .A(key[58]), .Y(n5477) );
  AOI221XL U3940 ( .A0(n1648), .A1(n22), .B0(n1630), .B1(key[186]), .C0(n5474), 
        .Y(n5475) );
  AO22X1 U3941 ( .A0(prev_key1_reg[58]), .A1(n1614), .B0(n1601), .B1(n5473), 
        .Y(n5474) );
  OAI221XL U3942 ( .A0(n1672), .A1(n5467), .B0(n5466), .B1(n1654), .C0(n5465), 
        .Y(n3822) );
  INVX1 U3943 ( .A(key[90]), .Y(n5467) );
  AOI221XL U3944 ( .A0(n1648), .A1(n895), .B0(n1630), .B1(key[218]), .C0(n5464), .Y(n5465) );
  AO22X1 U3945 ( .A0(prev_key1_reg[90]), .A1(n1614), .B0(n1601), .B1(n5463), 
        .Y(n5464) );
  OAI221XL U3946 ( .A0(n1671), .A1(n5418), .B0(n5417), .B1(n1656), .C0(n5416), 
        .Y(n3888) );
  INVX1 U3947 ( .A(key[24]), .Y(n5418) );
  AOI221XL U3948 ( .A0(n1645), .A1(n30), .B0(n1629), .B1(key[152]), .C0(n5415), 
        .Y(n5416) );
  AO22X1 U3949 ( .A0(sboxw[24]), .A1(n1613), .B0(n1600), .B1(n5414), .Y(n5415)
         );
  OAI221XL U3950 ( .A0(n1671), .A1(n5405), .B0(n5404), .B1(n1656), .C0(n5403), 
        .Y(n3856) );
  INVX1 U3951 ( .A(key[56]), .Y(n5405) );
  AOI221XL U3952 ( .A0(n1649), .A1(n23), .B0(n1629), .B1(key[184]), .C0(n5402), 
        .Y(n5403) );
  AO22X1 U3953 ( .A0(prev_key1_reg[56]), .A1(n1613), .B0(n1600), .B1(n5401), 
        .Y(n5402) );
  OAI221XL U3954 ( .A0(n1671), .A1(n5395), .B0(n5394), .B1(n1656), .C0(n5393), 
        .Y(n3824) );
  INVX1 U3955 ( .A(key[88]), .Y(n5395) );
  AOI221XL U3956 ( .A0(n1637), .A1(n903), .B0(n1629), .B1(key[216]), .C0(n5392), .Y(n5393) );
  AO22X1 U3957 ( .A0(prev_key1_reg[88]), .A1(n1613), .B0(n1600), .B1(n5391), 
        .Y(n5392) );
  OAI221XL U3958 ( .A0(n1664), .A1(n5648), .B0(n5647), .B1(n1654), .C0(n5646), 
        .Y(n3817) );
  INVX1 U3959 ( .A(key[95]), .Y(n5648) );
  INVX1 U3960 ( .A(n5683), .Y(n5647) );
  AOI221XL U3961 ( .A0(n1636), .A1(n5684), .B0(n1631), .B1(key[223]), .C0(
        n5645), .Y(n5646) );
  OAI221XL U3962 ( .A0(n1676), .A1(n5640), .B0(n1663), .B1(n5639), .C0(n5638), 
        .Y(n3785) );
  INVX1 U3963 ( .A(key[127]), .Y(n5640) );
  INVX1 U3964 ( .A(n5685), .Y(n5639) );
  AOI221XL U3965 ( .A0(n5686), .A1(n1636), .B0(n1635), .B1(key[255]), .C0(
        n5637), .Y(n5638) );
  OAI221XL U3966 ( .A0(n1664), .A1(n4761), .B0(n1659), .B1(n4760), .C0(n4759), 
        .Y(n3908) );
  INVX1 U3967 ( .A(key[4]), .Y(n4761) );
  INVX1 U3968 ( .A(n5742), .Y(n4760) );
  AOI221XL U3969 ( .A0(n1643), .A1(n36), .B0(n1623), .B1(key[132]), .C0(n4758), 
        .Y(n4759) );
  OAI221XL U3970 ( .A0(n1674), .A1(n5021), .B0(n1662), .B1(n5020), .C0(n5019), 
        .Y(n3900) );
  INVX1 U3971 ( .A(key[12]), .Y(n5021) );
  AOI221XL U3972 ( .A0(n1641), .A1(n33), .B0(n1625), .B1(key[140]), .C0(n5018), 
        .Y(n5019) );
  OAI221XL U3973 ( .A0(n1666), .A1(n4653), .B0(n1659), .B1(n4652), .C0(n4651), 
        .Y(n3879) );
  INVX1 U3974 ( .A(key[33]), .Y(n4653) );
  INVX1 U3975 ( .A(n5752), .Y(n4652) );
  AOI221XL U3976 ( .A0(n1646), .A1(n1123), .B0(n1622), .B1(key[161]), .C0(
        n4650), .Y(n4651) );
  OAI221XL U3977 ( .A0(n1664), .A1(n4685), .B0(n1660), .B1(n4684), .C0(n4683), 
        .Y(n3878) );
  INVX1 U3978 ( .A(key[34]), .Y(n4685) );
  INVX1 U3979 ( .A(n5749), .Y(n4684) );
  AOI221XL U3980 ( .A0(n1647), .A1(n1119), .B0(n1623), .B1(key[162]), .C0(
        n4682), .Y(n4683) );
  OAI221XL U3981 ( .A0(n1673), .A1(n4781), .B0(n1661), .B1(n4780), .C0(n4779), 
        .Y(n3875) );
  INVX1 U3982 ( .A(key[37]), .Y(n4781) );
  INVX1 U3983 ( .A(n5740), .Y(n4780) );
  AOI221XL U3984 ( .A0(n1643), .A1(n1107), .B0(n1624), .B1(key[165]), .C0(
        n4778), .Y(n4779) );
  OAI221XL U3985 ( .A0(n1667), .A1(n4844), .B0(n1660), .B1(n4843), .C0(n4842), 
        .Y(n3873) );
  INVX1 U3986 ( .A(key[39]), .Y(n4844) );
  INVX1 U3987 ( .A(n5734), .Y(n4843) );
  AOI221XL U3988 ( .A0(n1645), .A1(n1099), .B0(n1634), .B1(key[167]), .C0(
        n4841), .Y(n4842) );
  OAI221XL U3989 ( .A0(n1674), .A1(n5009), .B0(n1658), .B1(n5008), .C0(n5007), 
        .Y(n3868) );
  INVX1 U3990 ( .A(key[44]), .Y(n5009) );
  AOI221XL U3991 ( .A0(n1641), .A1(n1079), .B0(n1625), .B1(key[172]), .C0(
        n5006), .Y(n5007) );
  OAI221XL U3992 ( .A0(n1673), .A1(n5042), .B0(n1662), .B1(n5041), .C0(n5040), 
        .Y(n3867) );
  INVX1 U3993 ( .A(key[45]), .Y(n5042) );
  INVX1 U3994 ( .A(n5716), .Y(n5041) );
  AOI221XL U3995 ( .A0(n1641), .A1(n1075), .B0(n1625), .B1(key[173]), .C0(
        n5039), .Y(n5040) );
  OAI221XL U3996 ( .A0(n1670), .A1(n5272), .B0(n1651), .B1(n5271), .C0(n5270), 
        .Y(n3860) );
  INVX1 U3997 ( .A(key[52]), .Y(n5272) );
  AOI221XL U3998 ( .A0(n1638), .A1(n1047), .B0(n1628), .B1(key[180]), .C0(
        n5269), .Y(n5270) );
  OAI221XL U3999 ( .A0(n1667), .A1(n4902), .B0(n1661), .B1(n4901), .C0(n4900), 
        .Y(n3839) );
  INVX1 U4000 ( .A(key[73]), .Y(n4902) );
  AOI221XL U4001 ( .A0(n1648), .A1(n31), .B0(n1632), .B1(key[201]), .C0(n4899), 
        .Y(n4900) );
  OAI221XL U4002 ( .A0(n1670), .A1(n5264), .B0(n1651), .B1(n5263), .C0(n5262), 
        .Y(n3828) );
  INVX1 U4003 ( .A(key[84]), .Y(n5264) );
  AOI221XL U4004 ( .A0(n1638), .A1(n32), .B0(n1628), .B1(key[212]), .C0(n5261), 
        .Y(n5262) );
  INVX1 U4005 ( .A(n4951), .Y(n1213) );
  AOI222XL U4006 ( .A0(n1715), .A1(n55), .B0(key[10]), .B1(n1685), .C0(n1699), 
        .C1(n5724), .Y(n1214) );
  INVX1 U4007 ( .A(n5050), .Y(n1201) );
  AOI222XL U4008 ( .A0(n1716), .A1(n57), .B0(key[13]), .B1(n1685), .C0(n1699), 
        .C1(n5715), .Y(n1202) );
  INVX1 U4009 ( .A(n5214), .Y(n1181) );
  AOI222XL U4010 ( .A0(n1714), .A1(n58), .B0(key[18]), .B1(n1689), .C0(n1701), 
        .C1(n5701), .Y(n1182) );
  INVX1 U4011 ( .A(n4939), .Y(n1085) );
  AOI222XL U4012 ( .A0(n1711), .A1(n1087), .B0(key[42]), .B1(n1684), .C0(n1698), .C1(n5725), .Y(n1086) );
  INVX1 U4013 ( .A(n5038), .Y(n1073) );
  AOI222XL U4014 ( .A0(n1711), .A1(n1075), .B0(key[45]), .B1(n1684), .C0(n1698), .C1(n5716), .Y(n1074) );
  INVX1 U4015 ( .A(n5202), .Y(n1053) );
  AOI222XL U4016 ( .A0(n1710), .A1(n1055), .B0(key[50]), .B1(n1683), .C0(n1697), .C1(n5702), .Y(n1054) );
  INVX1 U4017 ( .A(n5301), .Y(n1041) );
  AOI222XL U4018 ( .A0(n1710), .A1(n1043), .B0(key[53]), .B1(n1683), .C0(n1697), .C1(n5693), .Y(n1042) );
  INVX1 U4019 ( .A(n5366), .Y(n1033) );
  AOI222XL U4020 ( .A0(n1710), .A1(n1035), .B0(key[55]), .B1(n1683), .C0(n1697), .C1(n5688), .Y(n1034) );
  INVX1 U4021 ( .A(n4931), .Y(n957) );
  AOI222XL U4022 ( .A0(n1708), .A1(n42), .B0(key[74]), .B1(n1690), .C0(n1695), 
        .C1(n5726), .Y(n958) );
  INVX1 U4023 ( .A(n5030), .Y(n945) );
  AOI222XL U4024 ( .A0(n1708), .A1(n44), .B0(key[77]), .B1(n1690), .C0(n1695), 
        .C1(n5717), .Y(n946) );
  INVX1 U4025 ( .A(n5095), .Y(n937) );
  AOI222XL U4026 ( .A0(n1707), .A1(n45), .B0(key[79]), .B1(n1682), .C0(n1703), 
        .C1(n5712), .Y(n938) );
  INVX1 U4027 ( .A(n5194), .Y(n925) );
  AOI222XL U4028 ( .A0(n1707), .A1(n46), .B0(key[82]), .B1(n1682), .C0(n1702), 
        .C1(n5703), .Y(n926) );
  INVX1 U4029 ( .A(n5293), .Y(n913) );
  AOI222XL U4030 ( .A0(n1707), .A1(n47), .B0(key[85]), .B1(n1682), .C0(n1697), 
        .C1(n5694), .Y(n914) );
  INVX1 U4031 ( .A(n5358), .Y(n905) );
  AOI222XL U4032 ( .A0(n1707), .A1(n48), .B0(key[87]), .B1(n1682), .C0(n1701), 
        .C1(n5689), .Y(n906) );
  AOI222XL U4033 ( .A0(n1705), .A1(n835), .B0(key[105]), .B1(n1680), .C0(n1693), .C1(n836), .Y(n834) );
  INVX1 U4034 ( .A(n4895), .Y(n836) );
  AOI222XL U4035 ( .A0(n1715), .A1(n5680), .B0(key[31]), .B1(n1688), .C0(n1699), .C1(n5679), .Y(n1130) );
  AOI222XL U4036 ( .A0(n1709), .A1(n5682), .B0(key[63]), .B1(n1686), .C0(n1696), .C1(n5681), .Y(n1002) );
  AOI222XL U4037 ( .A0(n1714), .A1(n16), .B0(key[1]), .B1(n1690), .C0(n1700), 
        .C1(n5751), .Y(n1250) );
  AOI222XL U4038 ( .A0(n1716), .A1(n36), .B0(key[4]), .B1(n1685), .C0(n1703), 
        .C1(n5742), .Y(n1238) );
  AOI222XL U4039 ( .A0(n1713), .A1(n1123), .B0(key[33]), .B1(n1687), .C0(n1700), .C1(n5752), .Y(n1122) );
  AOI222XL U4040 ( .A0(n1708), .A1(n1111), .B0(key[36]), .B1(n1686), .C0(n5758), .C1(n5743), .Y(n1110) );
  AOI222XL U4041 ( .A0(n1709), .A1(n15), .B0(key[65]), .B1(n5757), .C0(n1696), 
        .C1(n5753), .Y(n994) );
  AOI222XL U4042 ( .A0(n1709), .A1(n34), .B0(key[68]), .B1(n1683), .C0(n1696), 
        .C1(n5744), .Y(n982) );
  OAI221XL U4043 ( .A0(n1666), .A1(n4639), .B0(n4638), .B1(n1658), .C0(n4637), 
        .Y(n3815) );
  INVX1 U4044 ( .A(key[97]), .Y(n4639) );
  AOI221XL U4045 ( .A0(n1644), .A1(n867), .B0(n1622), .B1(key[225]), .C0(n4636), .Y(n4637) );
  OAI221XL U4046 ( .A0(n1666), .A1(n4671), .B0(n4670), .B1(n1658), .C0(n4669), 
        .Y(n3814) );
  INVX1 U4047 ( .A(key[98]), .Y(n4671) );
  AOI221XL U4048 ( .A0(n1644), .A1(n863), .B0(n1622), .B1(key[226]), .C0(n4668), .Y(n4669) );
  AO22X1 U4049 ( .A0(prev_key1_reg[98]), .A1(n1608), .B0(n1595), .B1(n4667), 
        .Y(n4668) );
  OAI221XL U4050 ( .A0(n1676), .A1(n4703), .B0(n4702), .B1(n1658), .C0(n4701), 
        .Y(n3813) );
  INVX1 U4051 ( .A(key[99]), .Y(n4703) );
  AOI221XL U4052 ( .A0(n1644), .A1(n859), .B0(n1623), .B1(key[227]), .C0(n4700), .Y(n4701) );
  AO22X1 U4053 ( .A0(prev_key1_reg[99]), .A1(n1618), .B0(n1606), .B1(n4699), 
        .Y(n4700) );
  OAI221XL U4054 ( .A0(n1677), .A1(n4735), .B0(n4734), .B1(n1658), .C0(n4733), 
        .Y(n3812) );
  INVX1 U4055 ( .A(key[100]), .Y(n4735) );
  AOI221XL U4056 ( .A0(n1644), .A1(n855), .B0(n1623), .B1(key[228]), .C0(n4732), .Y(n4733) );
  AO22X1 U4057 ( .A0(prev_key1_reg[100]), .A1(n1619), .B0(n1604), .B1(n4731), 
        .Y(n4732) );
  OAI221XL U4058 ( .A0(n1665), .A1(n4767), .B0(n4766), .B1(n1658), .C0(n4765), 
        .Y(n3811) );
  INVX1 U4059 ( .A(key[101]), .Y(n4767) );
  AOI221XL U4060 ( .A0(n1643), .A1(n851), .B0(n1624), .B1(key[229]), .C0(n4764), .Y(n4765) );
  AO22X1 U4061 ( .A0(prev_key1_reg[101]), .A1(n1620), .B0(n1606), .B1(n4763), 
        .Y(n4764) );
  OAI221XL U4062 ( .A0(n1665), .A1(n4830), .B0(n4829), .B1(n1658), .C0(n4828), 
        .Y(n3809) );
  INVX1 U4063 ( .A(key[103]), .Y(n4830) );
  AOI221XL U4064 ( .A0(n1643), .A1(n843), .B0(n1624), .B1(key[231]), .C0(n4827), .Y(n4828) );
  AO22X1 U4065 ( .A0(prev_key1_reg[103]), .A1(n1621), .B0(n1606), .B1(n4826), 
        .Y(n4827) );
  OAI221XL U4066 ( .A0(n1668), .A1(n4929), .B0(n4928), .B1(n1657), .C0(n4927), 
        .Y(n3806) );
  INVX1 U4067 ( .A(key[106]), .Y(n4929) );
  AOI221XL U4068 ( .A0(n1642), .A1(n831), .B0(n1634), .B1(key[234]), .C0(n4926), .Y(n4927) );
  AO22X1 U4069 ( .A0(prev_key1_reg[106]), .A1(n1619), .B0(n1604), .B1(n4925), 
        .Y(n4926) );
  OAI221XL U4070 ( .A0(n1677), .A1(n5028), .B0(n5027), .B1(n1657), .C0(n5026), 
        .Y(n3803) );
  INVX1 U4071 ( .A(key[109]), .Y(n5028) );
  AOI221XL U4072 ( .A0(n1641), .A1(n819), .B0(n1625), .B1(key[237]), .C0(n5025), .Y(n5026) );
  AO22X1 U4073 ( .A0(prev_key1_reg[109]), .A1(n1609), .B0(n1596), .B1(n5024), 
        .Y(n5025) );
  OAI221XL U4074 ( .A0(n1675), .A1(n5093), .B0(n5092), .B1(n1657), .C0(n5091), 
        .Y(n3801) );
  INVX1 U4075 ( .A(key[111]), .Y(n5093) );
  AOI221XL U4076 ( .A0(n1640), .A1(n811), .B0(n1626), .B1(key[239]), .C0(n5090), .Y(n5091) );
  AO22X1 U4077 ( .A0(prev_key1_reg[111]), .A1(n1610), .B0(n1597), .B1(n5089), 
        .Y(n5090) );
  OAI221XL U4078 ( .A0(n1675), .A1(n5126), .B0(n5125), .B1(n1657), .C0(n5124), 
        .Y(n3800) );
  INVX1 U4079 ( .A(key[112]), .Y(n5126) );
  AOI221XL U4080 ( .A0(n1640), .A1(n807), .B0(n1626), .B1(key[240]), .C0(n5123), .Y(n5124) );
  AO22X1 U4081 ( .A0(prev_key1_reg[112]), .A1(n1610), .B0(n1597), .B1(n5122), 
        .Y(n5123) );
  OAI221XL U4082 ( .A0(n1677), .A1(n5159), .B0(n5158), .B1(n1657), .C0(n5157), 
        .Y(n3799) );
  INVX1 U4083 ( .A(key[113]), .Y(n5159) );
  AOI221XL U4084 ( .A0(n1639), .A1(n803), .B0(n1626), .B1(key[241]), .C0(n5156), .Y(n5157) );
  AO22X1 U4085 ( .A0(prev_key1_reg[113]), .A1(n1610), .B0(n1597), .B1(n5155), 
        .Y(n5156) );
  OAI221XL U4086 ( .A0(n1669), .A1(n5192), .B0(n5191), .B1(n1657), .C0(n5190), 
        .Y(n3798) );
  INVX1 U4087 ( .A(key[114]), .Y(n5192) );
  AOI221XL U4088 ( .A0(n1639), .A1(n799), .B0(n1627), .B1(key[242]), .C0(n5189), .Y(n5190) );
  AO22X1 U4089 ( .A0(prev_key1_reg[114]), .A1(n1611), .B0(n1598), .B1(n5188), 
        .Y(n5189) );
  OAI221XL U4090 ( .A0(n1670), .A1(n5258), .B0(n5257), .B1(n1656), .C0(n5256), 
        .Y(n3796) );
  INVX1 U4091 ( .A(key[116]), .Y(n5258) );
  AOI221XL U4092 ( .A0(n1638), .A1(n791), .B0(n1628), .B1(key[244]), .C0(n5255), .Y(n5256) );
  AO22X1 U4093 ( .A0(prev_key1_reg[116]), .A1(n1612), .B0(n1599), .B1(n5254), 
        .Y(n5255) );
  OAI221XL U4094 ( .A0(n1670), .A1(n5291), .B0(n5290), .B1(n1656), .C0(n5289), 
        .Y(n3795) );
  INVX1 U4095 ( .A(key[117]), .Y(n5291) );
  AOI221XL U4096 ( .A0(n1638), .A1(n787), .B0(n1628), .B1(key[245]), .C0(n5288), .Y(n5289) );
  AO22X1 U4097 ( .A0(prev_key1_reg[117]), .A1(n1612), .B0(n1599), .B1(n5287), 
        .Y(n5288) );
  OAI221XL U4098 ( .A0(n1670), .A1(n5324), .B0(n5323), .B1(n1656), .C0(n5322), 
        .Y(n3794) );
  INVX1 U4099 ( .A(key[118]), .Y(n5324) );
  AOI221XL U4100 ( .A0(n1637), .A1(n783), .B0(n1628), .B1(key[246]), .C0(n5321), .Y(n5322) );
  AO22X1 U4101 ( .A0(prev_key1_reg[118]), .A1(n1612), .B0(n1599), .B1(n5320), 
        .Y(n5321) );
  OAI221XL U4102 ( .A0(n1671), .A1(n5356), .B0(n5355), .B1(n1656), .C0(n5354), 
        .Y(n3793) );
  INVX1 U4103 ( .A(key[119]), .Y(n5356) );
  AOI221XL U4104 ( .A0(n1637), .A1(n779), .B0(n1629), .B1(key[247]), .C0(n5353), .Y(n5354) );
  AO22X1 U4105 ( .A0(prev_key1_reg[119]), .A1(n1613), .B0(n1600), .B1(n5352), 
        .Y(n5353) );
  OAI221XL U4106 ( .A0(n1677), .A1(n5676), .B0(n5675), .B1(n1656), .C0(n5673), 
        .Y(n3881) );
  INVX1 U4107 ( .A(key[31]), .Y(n5676) );
  INVX1 U4108 ( .A(n5679), .Y(n5675) );
  AOI221XL U4109 ( .A0(n1640), .A1(n5680), .B0(n1632), .B1(key[159]), .C0(
        n5670), .Y(n5673) );
  OAI221XL U4110 ( .A0(n1675), .A1(n5657), .B0(n5656), .B1(n1655), .C0(n5655), 
        .Y(n3849) );
  INVX1 U4111 ( .A(key[63]), .Y(n5657) );
  INVX1 U4112 ( .A(n5681), .Y(n5656) );
  AOI221XL U4113 ( .A0(n1636), .A1(n5682), .B0(n1634), .B1(key[191]), .C0(
        n5654), .Y(n5655) );
  OAI221XL U4114 ( .A0(n1672), .A1(n5424), .B0(n5423), .B1(n1654), .C0(n5422), 
        .Y(n3791) );
  INVX1 U4115 ( .A(key[121]), .Y(n5424) );
  AOI221XL U4116 ( .A0(n1646), .A1(n59), .B0(n1630), .B1(key[249]), .C0(n5421), 
        .Y(n5422) );
  AO22X1 U4117 ( .A0(prev_key1_reg[121]), .A1(n1614), .B0(n1601), .B1(n5420), 
        .Y(n5421) );
  OAI221XL U4118 ( .A0(n1677), .A1(n5532), .B0(n5531), .B1(n1653), .C0(n5530), 
        .Y(n3788) );
  INVX1 U4119 ( .A(key[124]), .Y(n5532) );
  AOI221XL U4120 ( .A0(n1646), .A1(n60), .B0(n1633), .B1(key[252]), .C0(n5529), 
        .Y(n5530) );
  AO22X1 U4121 ( .A0(prev_key1_reg[124]), .A1(n1615), .B0(n1603), .B1(n5528), 
        .Y(n5529) );
  OAI221XL U4122 ( .A0(n1675), .A1(n5568), .B0(n5567), .B1(n1655), .C0(n5566), 
        .Y(n3787) );
  INVX1 U4123 ( .A(key[125]), .Y(n5568) );
  AOI221XL U4124 ( .A0(n1649), .A1(n61), .B0(n1632), .B1(key[253]), .C0(n5565), 
        .Y(n5566) );
  AO22X1 U4125 ( .A0(prev_key1_reg[125]), .A1(n1615), .B0(n5668), .B1(n5564), 
        .Y(n5565) );
  OAI221XL U4126 ( .A0(n1664), .A1(n5604), .B0(n5603), .B1(n1654), .C0(n5602), 
        .Y(n3786) );
  INVX1 U4127 ( .A(key[126]), .Y(n5604) );
  AOI221XL U4128 ( .A0(n1636), .A1(n62), .B0(n1631), .B1(key[254]), .C0(n5601), 
        .Y(n5602) );
  AO22X1 U4129 ( .A0(prev_key1_reg[126]), .A1(n1616), .B0(n1602), .B1(n5600), 
        .Y(n5601) );
  OAI221XL U4130 ( .A0(n1672), .A1(n5496), .B0(n5495), .B1(n1654), .C0(n5494), 
        .Y(n3789) );
  INVX1 U4131 ( .A(key[123]), .Y(n5496) );
  AOI221XL U4132 ( .A0(n1647), .A1(n63), .B0(n1630), .B1(key[251]), .C0(n5493), 
        .Y(n5494) );
  AO22X1 U4133 ( .A0(prev_key1_reg[123]), .A1(n1614), .B0(n1601), .B1(n5492), 
        .Y(n5493) );
  OAI221XL U4134 ( .A0(n1672), .A1(n5460), .B0(n5459), .B1(n1655), .C0(n5458), 
        .Y(n3790) );
  INVX1 U4135 ( .A(key[122]), .Y(n5460) );
  AOI221XL U4136 ( .A0(n5672), .A1(n64), .B0(n1630), .B1(key[250]), .C0(n5457), 
        .Y(n5458) );
  AO22X1 U4137 ( .A0(prev_key1_reg[122]), .A1(n1614), .B0(n1601), .B1(n5456), 
        .Y(n5457) );
  OAI221XL U4138 ( .A0(n1671), .A1(n5388), .B0(n5387), .B1(n1656), .C0(n5386), 
        .Y(n3792) );
  INVX1 U4139 ( .A(key[120]), .Y(n5388) );
  AOI221XL U4140 ( .A0(n1637), .A1(n65), .B0(n1629), .B1(key[248]), .C0(n5385), 
        .Y(n5386) );
  AO22X1 U4141 ( .A0(prev_key1_reg[120]), .A1(n1613), .B0(n1600), .B1(n5384), 
        .Y(n5385) );
  OAI221XL U4142 ( .A0(n1666), .A1(n4665), .B0(n1660), .B1(n4664), .C0(n4663), 
        .Y(n3911) );
  INVX1 U4143 ( .A(key[1]), .Y(n4665) );
  INVX1 U4144 ( .A(n5751), .Y(n4664) );
  AOI221XL U4145 ( .A0(n1645), .A1(n16), .B0(n1622), .B1(key[129]), .C0(n4662), 
        .Y(n4663) );
  OAI221XL U4146 ( .A0(n1665), .A1(n4697), .B0(n1653), .B1(n4696), .C0(n4695), 
        .Y(n3910) );
  INVX1 U4147 ( .A(key[2]), .Y(n4697) );
  INVX1 U4148 ( .A(n5748), .Y(n4696) );
  AOI221XL U4149 ( .A0(n1644), .A1(n50), .B0(n1623), .B1(key[130]), .C0(n4694), 
        .Y(n4695) );
  OAI221XL U4150 ( .A0(n1673), .A1(n4729), .B0(n1661), .B1(n4728), .C0(n4727), 
        .Y(n3909) );
  INVX1 U4151 ( .A(key[3]), .Y(n4729) );
  INVX1 U4152 ( .A(n5745), .Y(n4728) );
  AOI221XL U4153 ( .A0(n1644), .A1(n51), .B0(n1623), .B1(key[131]), .C0(n4726), 
        .Y(n4727) );
  OAI221XL U4154 ( .A0(n1664), .A1(n4793), .B0(n1661), .B1(n4792), .C0(n4791), 
        .Y(n3907) );
  INVX1 U4155 ( .A(key[5]), .Y(n4793) );
  INVX1 U4156 ( .A(n5739), .Y(n4792) );
  AOI221XL U4157 ( .A0(n1643), .A1(n52), .B0(n1624), .B1(key[133]), .C0(n4790), 
        .Y(n4791) );
  OAI221XL U4158 ( .A0(n1667), .A1(n4856), .B0(n1663), .B1(n4855), .C0(n4854), 
        .Y(n3905) );
  INVX1 U4159 ( .A(key[7]), .Y(n4856) );
  INVX1 U4160 ( .A(n5733), .Y(n4855) );
  AOI221XL U4161 ( .A0(n1646), .A1(n54), .B0(n1635), .B1(key[135]), .C0(n4853), 
        .Y(n4854) );
  OAI221XL U4162 ( .A0(n1667), .A1(n4922), .B0(n1663), .B1(n4921), .C0(n4920), 
        .Y(n3903) );
  INVX1 U4163 ( .A(key[9]), .Y(n4922) );
  AOI221XL U4164 ( .A0(n1642), .A1(n70), .B0(n1631), .B1(key[137]), .C0(n4919), 
        .Y(n4920) );
  OAI221XL U4165 ( .A0(n1668), .A1(n4955), .B0(n1663), .B1(n4954), .C0(n4953), 
        .Y(n3902) );
  INVX1 U4166 ( .A(key[10]), .Y(n4955) );
  INVX1 U4167 ( .A(n5724), .Y(n4954) );
  AOI221XL U4168 ( .A0(n1642), .A1(n55), .B0(n1634), .B1(key[138]), .C0(n4952), 
        .Y(n4953) );
  OAI221XL U4169 ( .A0(n1673), .A1(n5054), .B0(n1658), .B1(n5053), .C0(n5052), 
        .Y(n3899) );
  INVX1 U4170 ( .A(key[13]), .Y(n5054) );
  INVX1 U4171 ( .A(n5715), .Y(n5053) );
  AOI221XL U4172 ( .A0(n1641), .A1(n57), .B0(n1625), .B1(key[141]), .C0(n5051), 
        .Y(n5052) );
  OAI221XL U4173 ( .A0(n1676), .A1(n5119), .B0(n1652), .B1(n5118), .C0(n5117), 
        .Y(n3897) );
  INVX1 U4174 ( .A(key[15]), .Y(n5119) );
  INVX1 U4175 ( .A(n5710), .Y(n5118) );
  AOI221XL U4176 ( .A0(n1640), .A1(n12), .B0(n1626), .B1(key[143]), .C0(n5116), 
        .Y(n5117) );
  OAI221XL U4177 ( .A0(n1675), .A1(n5152), .B0(n1652), .B1(n5151), .C0(n5150), 
        .Y(n3896) );
  INVX1 U4178 ( .A(key[16]), .Y(n5152) );
  AOI221XL U4179 ( .A0(n1640), .A1(n71), .B0(n1626), .B1(key[144]), .C0(n5149), 
        .Y(n5150) );
  OAI221XL U4180 ( .A0(n1669), .A1(n5185), .B0(n1651), .B1(n5184), .C0(n5183), 
        .Y(n3895) );
  INVX1 U4181 ( .A(key[17]), .Y(n5185) );
  INVX1 U4182 ( .A(n5704), .Y(n5184) );
  AOI221XL U4183 ( .A0(n1639), .A1(n72), .B0(n1627), .B1(key[145]), .C0(n5182), 
        .Y(n5183) );
  OAI221XL U4184 ( .A0(n1669), .A1(n5218), .B0(n1651), .B1(n5217), .C0(n5216), 
        .Y(n3894) );
  INVX1 U4185 ( .A(key[18]), .Y(n5218) );
  INVX1 U4186 ( .A(n5701), .Y(n5217) );
  AOI221XL U4187 ( .A0(n1639), .A1(n58), .B0(n1627), .B1(key[146]), .C0(n5215), 
        .Y(n5216) );
  OAI221XL U4188 ( .A0(n1670), .A1(n5284), .B0(n1650), .B1(n5283), .C0(n5282), 
        .Y(n3892) );
  INVX1 U4189 ( .A(key[20]), .Y(n5284) );
  AOI221XL U4190 ( .A0(n1638), .A1(n73), .B0(n1628), .B1(key[148]), .C0(n5281), 
        .Y(n5282) );
  OAI221XL U4191 ( .A0(n1670), .A1(n5317), .B0(n1650), .B1(n5316), .C0(n5315), 
        .Y(n3891) );
  INVX1 U4192 ( .A(key[21]), .Y(n5317) );
  INVX1 U4193 ( .A(n5692), .Y(n5316) );
  AOI221XL U4194 ( .A0(n1638), .A1(n13), .B0(n1628), .B1(key[149]), .C0(n5314), 
        .Y(n5315) );
  OAI221XL U4195 ( .A0(n1671), .A1(n5349), .B0(n1650), .B1(n5348), .C0(n5347), 
        .Y(n3890) );
  INVX1 U4196 ( .A(key[22]), .Y(n5349) );
  AOI221XL U4197 ( .A0(n1637), .A1(n74), .B0(n1629), .B1(key[150]), .C0(n5346), 
        .Y(n5347) );
  OAI221XL U4198 ( .A0(n1671), .A1(n5382), .B0(n1650), .B1(n5381), .C0(n5380), 
        .Y(n3889) );
  INVX1 U4199 ( .A(key[23]), .Y(n5382) );
  INVX1 U4200 ( .A(n5687), .Y(n5381) );
  AOI221XL U4201 ( .A0(n1637), .A1(n14), .B0(n1629), .B1(key[151]), .C0(n5379), 
        .Y(n5380) );
  OAI221XL U4202 ( .A0(n1666), .A1(n4645), .B0(n1653), .B1(n4644), .C0(n4643), 
        .Y(n3847) );
  INVX1 U4203 ( .A(key[65]), .Y(n4645) );
  INVX1 U4204 ( .A(n5753), .Y(n4644) );
  AOI221XL U4205 ( .A0(n1649), .A1(n15), .B0(n1622), .B1(key[193]), .C0(n4642), 
        .Y(n4643) );
  OAI221XL U4206 ( .A0(n1666), .A1(n4677), .B0(n1663), .B1(n4676), .C0(n4675), 
        .Y(n3846) );
  INVX1 U4207 ( .A(key[66]), .Y(n4677) );
  INVX1 U4208 ( .A(n5750), .Y(n4676) );
  AOI221XL U4209 ( .A0(n1644), .A1(n37), .B0(n1622), .B1(key[194]), .C0(n4674), 
        .Y(n4675) );
  OAI221XL U4210 ( .A0(n1674), .A1(n4709), .B0(n1660), .B1(n4708), .C0(n4707), 
        .Y(n3845) );
  INVX1 U4211 ( .A(key[67]), .Y(n4709) );
  INVX1 U4212 ( .A(n5747), .Y(n4708) );
  AOI221XL U4213 ( .A0(n1644), .A1(n38), .B0(n1623), .B1(key[195]), .C0(n4706), 
        .Y(n4707) );
  OAI221XL U4214 ( .A0(n1674), .A1(n4773), .B0(n1662), .B1(n4772), .C0(n4771), 
        .Y(n3843) );
  INVX1 U4215 ( .A(key[69]), .Y(n4773) );
  INVX1 U4216 ( .A(n5741), .Y(n4772) );
  AOI221XL U4217 ( .A0(n1643), .A1(n39), .B0(n1624), .B1(key[197]), .C0(n4770), 
        .Y(n4771) );
  OAI221XL U4218 ( .A0(n1665), .A1(n4836), .B0(n1661), .B1(n4835), .C0(n4834), 
        .Y(n3841) );
  INVX1 U4219 ( .A(key[71]), .Y(n4836) );
  INVX1 U4220 ( .A(n5735), .Y(n4835) );
  AOI221XL U4221 ( .A0(n1644), .A1(n41), .B0(n1624), .B1(key[199]), .C0(n4833), 
        .Y(n4834) );
  OAI221XL U4222 ( .A0(n1668), .A1(n4935), .B0(n1660), .B1(n4934), .C0(n4933), 
        .Y(n3838) );
  INVX1 U4223 ( .A(key[74]), .Y(n4935) );
  INVX1 U4224 ( .A(n5726), .Y(n4934) );
  AOI221XL U4225 ( .A0(n1642), .A1(n42), .B0(n1633), .B1(key[202]), .C0(n4932), 
        .Y(n4933) );
  OAI221XL U4226 ( .A0(n1668), .A1(n5001), .B0(n1661), .B1(n5000), .C0(n4999), 
        .Y(n3836) );
  INVX1 U4227 ( .A(key[76]), .Y(n5001) );
  AOI221XL U4228 ( .A0(n1641), .A1(n69), .B0(n1632), .B1(key[204]), .C0(n4998), 
        .Y(n4999) );
  OAI221XL U4229 ( .A0(n1677), .A1(n5034), .B0(n1659), .B1(n5033), .C0(n5032), 
        .Y(n3835) );
  INVX1 U4230 ( .A(key[77]), .Y(n5034) );
  INVX1 U4231 ( .A(n5717), .Y(n5033) );
  AOI221XL U4232 ( .A0(n1641), .A1(n44), .B0(n1625), .B1(key[205]), .C0(n5031), 
        .Y(n5032) );
  OAI221XL U4233 ( .A0(n1677), .A1(n5099), .B0(n1652), .B1(n5098), .C0(n5097), 
        .Y(n3833) );
  INVX1 U4234 ( .A(key[79]), .Y(n5099) );
  INVX1 U4235 ( .A(n5712), .Y(n5098) );
  AOI221XL U4236 ( .A0(n1640), .A1(n45), .B0(n1626), .B1(key[207]), .C0(n5096), 
        .Y(n5097) );
  OAI221XL U4237 ( .A0(n1676), .A1(n5132), .B0(n1652), .B1(n5131), .C0(n5130), 
        .Y(n3832) );
  INVX1 U4238 ( .A(key[80]), .Y(n5132) );
  AOI221XL U4239 ( .A0(n1640), .A1(n66), .B0(n1626), .B1(key[208]), .C0(n5129), 
        .Y(n5130) );
  OAI221XL U4240 ( .A0(n1674), .A1(n5165), .B0(n1652), .B1(n5164), .C0(n5163), 
        .Y(n3831) );
  INVX1 U4241 ( .A(key[81]), .Y(n5165) );
  INVX1 U4242 ( .A(n5706), .Y(n5164) );
  AOI221XL U4243 ( .A0(n1639), .A1(n67), .B0(n1626), .B1(key[209]), .C0(n5162), 
        .Y(n5163) );
  OAI221XL U4244 ( .A0(n1669), .A1(n5198), .B0(n1651), .B1(n5197), .C0(n5196), 
        .Y(n3830) );
  INVX1 U4245 ( .A(key[82]), .Y(n5198) );
  INVX1 U4246 ( .A(n5703), .Y(n5197) );
  AOI221XL U4247 ( .A0(n1639), .A1(n46), .B0(n1627), .B1(key[210]), .C0(n5195), 
        .Y(n5196) );
  OAI221XL U4248 ( .A0(n1670), .A1(n5297), .B0(n1650), .B1(n5296), .C0(n5295), 
        .Y(n3827) );
  INVX1 U4249 ( .A(key[85]), .Y(n5297) );
  INVX1 U4250 ( .A(n5694), .Y(n5296) );
  AOI221XL U4251 ( .A0(n1638), .A1(n47), .B0(n1628), .B1(key[213]), .C0(n5294), 
        .Y(n5295) );
  OAI221XL U4252 ( .A0(n1670), .A1(n5330), .B0(n1650), .B1(n5329), .C0(n5328), 
        .Y(n3826) );
  INVX1 U4253 ( .A(key[86]), .Y(n5330) );
  INVX1 U4254 ( .A(n5691), .Y(n5329) );
  AOI221XL U4255 ( .A0(n1637), .A1(n68), .B0(n1628), .B1(key[214]), .C0(n5327), 
        .Y(n5328) );
  OAI221XL U4256 ( .A0(n1671), .A1(n5362), .B0(n1650), .B1(n5361), .C0(n5360), 
        .Y(n3825) );
  INVX1 U4257 ( .A(key[87]), .Y(n5362) );
  INVX1 U4258 ( .A(n5689), .Y(n5361) );
  AOI221XL U4259 ( .A0(n1637), .A1(n48), .B0(n1629), .B1(key[215]), .C0(n5359), 
        .Y(n5360) );
  OAI221XL U4260 ( .A0(n1674), .A1(n4717), .B0(n1659), .B1(n4716), .C0(n4715), 
        .Y(n3877) );
  INVX1 U4261 ( .A(key[35]), .Y(n4717) );
  INVX1 U4262 ( .A(n5746), .Y(n4716) );
  AOI221XL U4263 ( .A0(n1645), .A1(n1115), .B0(n1623), .B1(key[163]), .C0(
        n4714), .Y(n4715) );
  OAI221XL U4264 ( .A0(n1673), .A1(n4749), .B0(n1662), .B1(n4748), .C0(n4747), 
        .Y(n3876) );
  INVX1 U4265 ( .A(key[36]), .Y(n4749) );
  INVX1 U4266 ( .A(n5743), .Y(n4748) );
  AOI221XL U4267 ( .A0(n1646), .A1(n1111), .B0(n1623), .B1(key[164]), .C0(
        n4746), .Y(n4747) );
  OAI221XL U4268 ( .A0(n1667), .A1(n4910), .B0(n1659), .B1(n4909), .C0(n4908), 
        .Y(n3871) );
  INVX1 U4269 ( .A(key[41]), .Y(n4910) );
  AOI221XL U4270 ( .A0(n1649), .A1(n1091), .B0(n1632), .B1(key[169]), .C0(
        n4907), .Y(n4908) );
  OAI221XL U4271 ( .A0(n1668), .A1(n4943), .B0(n1663), .B1(n4942), .C0(n4941), 
        .Y(n3870) );
  INVX1 U4272 ( .A(key[42]), .Y(n4943) );
  INVX1 U4273 ( .A(n5725), .Y(n4942) );
  AOI221XL U4274 ( .A0(n1642), .A1(n1087), .B0(n5671), .B1(key[170]), .C0(
        n4940), .Y(n4941) );
  OAI221XL U4275 ( .A0(n1673), .A1(n5107), .B0(n1652), .B1(n5106), .C0(n5105), 
        .Y(n3865) );
  INVX1 U4276 ( .A(key[47]), .Y(n5107) );
  INVX1 U4277 ( .A(n5711), .Y(n5106) );
  AOI221XL U4278 ( .A0(n1640), .A1(n1067), .B0(n1626), .B1(key[175]), .C0(
        n5104), .Y(n5105) );
  OAI221XL U4279 ( .A0(n1675), .A1(n5140), .B0(n1652), .B1(n5139), .C0(n5138), 
        .Y(n3864) );
  INVX1 U4280 ( .A(key[48]), .Y(n5140) );
  AOI221XL U4281 ( .A0(n1640), .A1(n1063), .B0(n1626), .B1(key[176]), .C0(
        n5137), .Y(n5138) );
  OAI221XL U4282 ( .A0(n1669), .A1(n5173), .B0(n1651), .B1(n5172), .C0(n5171), 
        .Y(n3863) );
  INVX1 U4283 ( .A(key[49]), .Y(n5173) );
  AOI221XL U4284 ( .A0(n1639), .A1(n1059), .B0(n1627), .B1(key[177]), .C0(
        n5170), .Y(n5171) );
  OAI221XL U4285 ( .A0(n1669), .A1(n5206), .B0(n1651), .B1(n5205), .C0(n5204), 
        .Y(n3862) );
  INVX1 U4286 ( .A(key[50]), .Y(n5206) );
  INVX1 U4287 ( .A(n5702), .Y(n5205) );
  AOI221XL U4288 ( .A0(n1639), .A1(n1055), .B0(n1627), .B1(key[178]), .C0(
        n5203), .Y(n5204) );
  OAI221XL U4289 ( .A0(n1670), .A1(n5305), .B0(n1650), .B1(n5304), .C0(n5303), 
        .Y(n3859) );
  INVX1 U4290 ( .A(key[53]), .Y(n5305) );
  INVX1 U4291 ( .A(n5693), .Y(n5304) );
  AOI221XL U4292 ( .A0(n1638), .A1(n1043), .B0(n1628), .B1(key[181]), .C0(
        n5302), .Y(n5303) );
  OAI221XL U4293 ( .A0(n1671), .A1(n5370), .B0(n1650), .B1(n5369), .C0(n5368), 
        .Y(n3857) );
  INVX1 U4294 ( .A(key[55]), .Y(n5370) );
  INVX1 U4295 ( .A(n5688), .Y(n5369) );
  AOI221XL U4296 ( .A0(n1637), .A1(n1035), .B0(n1629), .B1(key[183]), .C0(
        n5367), .Y(n5368) );
  OAI221XL U4297 ( .A0(n1671), .A1(n5337), .B0(n1650), .B1(n5), .C0(n5336), 
        .Y(n3858) );
  AOI221XL U4298 ( .A0(n1637), .A1(n1039), .B0(n1629), .B1(key[182]), .C0(
        n5335), .Y(n5336) );
  AO22X1 U4299 ( .A0(prev_key1_reg[54]), .A1(n1613), .B0(n1600), .B1(n5334), 
        .Y(n5335) );
  INVX1 U4300 ( .A(n5342), .Y(n1039) );
  XOR2X1 U4301 ( .A(n5419), .B(prev_key0_reg[121]), .Y(n769) );
  XOR2X1 U4302 ( .A(n5527), .B(prev_key0_reg[124]), .Y(n757) );
  XOR2X1 U4303 ( .A(n5563), .B(prev_key0_reg[125]), .Y(n753) );
  XOR2X1 U4304 ( .A(n5599), .B(prev_key0_reg[126]), .Y(n749) );
  XOR2X1 U4305 ( .A(n5491), .B(prev_key0_reg[123]), .Y(n761) );
  XOR2X1 U4306 ( .A(n5455), .B(prev_key0_reg[122]), .Y(n765) );
  XOR2X1 U4307 ( .A(n5383), .B(prev_key0_reg[120]), .Y(n773) );
  XOR2X1 U4308 ( .A(n5455), .B(prev_key0_reg[98]), .Y(n4670) );
  OAI221XL U4309 ( .A0(n1673), .A1(n4741), .B0(n1663), .B1(n4740), .C0(n4739), 
        .Y(n3844) );
  INVX1 U4310 ( .A(key[68]), .Y(n4741) );
  INVX1 U4311 ( .A(n5744), .Y(n4740) );
  AOI221XL U4312 ( .A0(n1645), .A1(n34), .B0(n1623), .B1(key[196]), .C0(n4738), 
        .Y(n4739) );
  AO22X1 U4313 ( .A0(prev_key1_reg[68]), .A1(n1617), .B0(n1606), .B1(n4737), 
        .Y(n4738) );
  OAI222XL U4314 ( .A0(n5884), .A1(n1589), .B0(n5662), .B1(n1572), .C0(n1566), 
        .C1(n5660), .Y(n3753) );
  INVX1 U4315 ( .A(prev_key0_reg[31]), .Y(n5660) );
  INVX1 U4316 ( .A(sboxw[31]), .Y(n5662) );
  OAI222XL U4317 ( .A0(n5771), .A1(n1587), .B0(n1574), .B1(n5445), .C0(n1555), 
        .C1(n5444), .Y(n3759) );
  INVX1 U4318 ( .A(prev_key0_reg[25]), .Y(n5444) );
  INVX1 U4319 ( .A(sboxw[25]), .Y(n5445) );
  OAI222XL U4320 ( .A0(n5769), .A1(n1587), .B0(n1575), .B1(n5443), .C0(n1555), 
        .C1(n5442), .Y(n3727) );
  INVX1 U4321 ( .A(prev_key0_reg[57]), .Y(n5442) );
  INVX1 U4322 ( .A(prev_key1_reg[57]), .Y(n5443) );
  OAI222XL U4323 ( .A0(n5770), .A1(n1587), .B0(n1574), .B1(n5433), .C0(n1555), 
        .C1(n5432), .Y(n3695) );
  INVX1 U4324 ( .A(prev_key0_reg[89]), .Y(n5432) );
  INVX1 U4325 ( .A(prev_key1_reg[89]), .Y(n5433) );
  OAI222XL U4326 ( .A0(n5836), .A1(n1588), .B0(n1573), .B1(n5553), .C0(n1554), 
        .C1(n5552), .Y(n3756) );
  INVX1 U4327 ( .A(prev_key0_reg[28]), .Y(n5552) );
  INVX1 U4328 ( .A(sboxw[28]), .Y(n5553) );
  OAI222XL U4329 ( .A0(n5834), .A1(n1588), .B0(n1573), .B1(n5551), .C0(n1554), 
        .C1(n5550), .Y(n3724) );
  INVX1 U4330 ( .A(prev_key0_reg[60]), .Y(n5550) );
  INVX1 U4331 ( .A(prev_key1_reg[60]), .Y(n5551) );
  OAI222XL U4332 ( .A0(n5832), .A1(n1588), .B0(n1573), .B1(n5541), .C0(n1554), 
        .C1(n5540), .Y(n3692) );
  INVX1 U4333 ( .A(prev_key0_reg[92]), .Y(n5540) );
  INVX1 U4334 ( .A(prev_key1_reg[92]), .Y(n5541) );
  OAI222XL U4335 ( .A0(n5852), .A1(n1588), .B0(n1572), .B1(n5589), .C0(n1553), 
        .C1(n5588), .Y(n3755) );
  INVX1 U4336 ( .A(prev_key0_reg[29]), .Y(n5588) );
  INVX1 U4337 ( .A(sboxw[29]), .Y(n5589) );
  OAI222XL U4338 ( .A0(n5850), .A1(n1588), .B0(n1573), .B1(n5587), .C0(n1553), 
        .C1(n5586), .Y(n3723) );
  INVX1 U4339 ( .A(prev_key0_reg[61]), .Y(n5586) );
  INVX1 U4340 ( .A(prev_key1_reg[61]), .Y(n5587) );
  OAI222XL U4341 ( .A0(n5848), .A1(n1588), .B0(n1573), .B1(n5577), .C0(n1554), 
        .C1(n5576), .Y(n3691) );
  INVX1 U4342 ( .A(prev_key0_reg[93]), .Y(n5576) );
  INVX1 U4343 ( .A(prev_key1_reg[93]), .Y(n5577) );
  OAI222XL U4344 ( .A0(n5868), .A1(n1589), .B0(n1573), .B1(n5625), .C0(n1553), 
        .C1(n5624), .Y(n3754) );
  INVX1 U4345 ( .A(prev_key0_reg[30]), .Y(n5624) );
  INVX1 U4346 ( .A(sboxw[30]), .Y(n5625) );
  OAI222XL U4347 ( .A0(n5866), .A1(n1589), .B0(n1572), .B1(n5623), .C0(n1553), 
        .C1(n5622), .Y(n3722) );
  INVX1 U4348 ( .A(prev_key0_reg[62]), .Y(n5622) );
  INVX1 U4349 ( .A(prev_key1_reg[62]), .Y(n5623) );
  OAI222XL U4350 ( .A0(n5864), .A1(n1589), .B0(n1575), .B1(n5613), .C0(n1553), 
        .C1(n5612), .Y(n3690) );
  INVX1 U4351 ( .A(prev_key0_reg[94]), .Y(n5612) );
  INVX1 U4352 ( .A(prev_key1_reg[94]), .Y(n5613) );
  OAI222XL U4353 ( .A0(n5820), .A1(n1588), .B0(n1574), .B1(n5517), .C0(n1554), 
        .C1(n5516), .Y(n3757) );
  INVX1 U4354 ( .A(prev_key0_reg[27]), .Y(n5516) );
  INVX1 U4355 ( .A(sboxw[27]), .Y(n5517) );
  OAI222XL U4356 ( .A0(n5818), .A1(n1588), .B0(n1573), .B1(n5515), .C0(n1554), 
        .C1(n5514), .Y(n3725) );
  INVX1 U4357 ( .A(prev_key0_reg[59]), .Y(n5514) );
  INVX1 U4358 ( .A(prev_key1_reg[59]), .Y(n5515) );
  OAI222XL U4359 ( .A0(n5816), .A1(n1587), .B0(n1574), .B1(n5505), .C0(n1554), 
        .C1(n5504), .Y(n3693) );
  INVX1 U4360 ( .A(prev_key0_reg[91]), .Y(n5504) );
  INVX1 U4361 ( .A(prev_key1_reg[91]), .Y(n5505) );
  OAI222XL U4362 ( .A0(n5804), .A1(n1587), .B0(n1574), .B1(n5481), .C0(n1555), 
        .C1(n5480), .Y(n3758) );
  INVX1 U4363 ( .A(prev_key0_reg[26]), .Y(n5480) );
  INVX1 U4364 ( .A(sboxw[26]), .Y(n5481) );
  OAI222XL U4365 ( .A0(n5802), .A1(n1587), .B0(n1574), .B1(n5479), .C0(n1555), 
        .C1(n5478), .Y(n3726) );
  INVX1 U4366 ( .A(prev_key0_reg[58]), .Y(n5478) );
  INVX1 U4367 ( .A(prev_key1_reg[58]), .Y(n5479) );
  OAI222XL U4368 ( .A0(n5800), .A1(n1587), .B0(n1574), .B1(n5469), .C0(n1555), 
        .C1(n5468), .Y(n3694) );
  INVX1 U4369 ( .A(prev_key0_reg[90]), .Y(n5468) );
  INVX1 U4370 ( .A(prev_key1_reg[90]), .Y(n5469) );
  OAI222XL U4371 ( .A0(n5788), .A1(n1586), .B0(n1575), .B1(n5409), .C0(n1555), 
        .C1(n5408), .Y(n3760) );
  INVX1 U4372 ( .A(prev_key0_reg[24]), .Y(n5408) );
  INVX1 U4373 ( .A(sboxw[24]), .Y(n5409) );
  OAI222XL U4374 ( .A0(n5786), .A1(n1586), .B0(n1575), .B1(n5407), .C0(n1555), 
        .C1(n5406), .Y(n3728) );
  INVX1 U4375 ( .A(prev_key0_reg[56]), .Y(n5406) );
  INVX1 U4376 ( .A(prev_key1_reg[56]), .Y(n5407) );
  OAI222XL U4377 ( .A0(n5784), .A1(n1586), .B0(n1569), .B1(n5397), .C0(n1563), 
        .C1(n5396), .Y(n3696) );
  INVX1 U4378 ( .A(prev_key0_reg[88]), .Y(n5396) );
  INVX1 U4379 ( .A(prev_key1_reg[88]), .Y(n5397) );
  OAI222XL U4380 ( .A0(n5882), .A1(n1589), .B0(n1572), .B1(n5659), .C0(n1553), 
        .C1(n5658), .Y(n3721) );
  INVX1 U4381 ( .A(prev_key0_reg[63]), .Y(n5658) );
  INVX1 U4382 ( .A(prev_key1_reg[63]), .Y(n5659) );
  OAI222XL U4383 ( .A0(n5880), .A1(n1589), .B0(n1572), .B1(n5650), .C0(n1553), 
        .C1(n5649), .Y(n3689) );
  INVX1 U4384 ( .A(prev_key0_reg[95]), .Y(n5649) );
  INVX1 U4385 ( .A(prev_key1_reg[95]), .Y(n5650) );
  OAI222XL U4386 ( .A0(n5790), .A1(n1581), .B0(n1567), .B1(n4625), .C0(n1565), 
        .C1(n4624), .Y(n3784) );
  INVX1 U4387 ( .A(prev_key0_reg[0]), .Y(n4624) );
  INVX1 U4388 ( .A(sboxw[0]), .Y(n4625) );
  OAI222XL U4389 ( .A0(n5781), .A1(n1581), .B0(n1577), .B1(n4657), .C0(n1566), 
        .C1(n4656), .Y(n3783) );
  INVX1 U4390 ( .A(prev_key0_reg[1]), .Y(n4656) );
  INVX1 U4391 ( .A(sboxw[1]), .Y(n4657) );
  OAI222XL U4392 ( .A0(n5806), .A1(n1590), .B0(n1567), .B1(n4689), .C0(n1557), 
        .C1(n4688), .Y(n3782) );
  INVX1 U4393 ( .A(prev_key0_reg[2]), .Y(n4688) );
  INVX1 U4394 ( .A(sboxw[2]), .Y(n4689) );
  OAI222XL U4395 ( .A0(n5822), .A1(n1592), .B0(n1567), .B1(n4721), .C0(n1565), 
        .C1(n4720), .Y(n3781) );
  INVX1 U4396 ( .A(prev_key0_reg[3]), .Y(n4720) );
  INVX1 U4397 ( .A(sboxw[3]), .Y(n4721) );
  OAI222XL U4398 ( .A0(n5838), .A1(n1591), .B0(n1579), .B1(n4753), .C0(n1566), 
        .C1(n4752), .Y(n3780) );
  INVX1 U4399 ( .A(prev_key0_reg[4]), .Y(n4752) );
  INVX1 U4400 ( .A(sboxw[4]), .Y(n4753) );
  OAI222XL U4401 ( .A0(n5854), .A1(n1591), .B0(n1568), .B1(n4785), .C0(n1557), 
        .C1(n4784), .Y(n3779) );
  INVX1 U4402 ( .A(prev_key0_reg[5]), .Y(n4784) );
  INVX1 U4403 ( .A(sboxw[5]), .Y(n4785) );
  OAI222XL U4404 ( .A0(n5870), .A1(n1594), .B0(n1567), .B1(n4816), .C0(n1557), 
        .C1(n4815), .Y(n3778) );
  INVX1 U4405 ( .A(prev_key0_reg[6]), .Y(n4815) );
  INVX1 U4406 ( .A(sboxw[6]), .Y(n4816) );
  OAI222XL U4407 ( .A0(n5886), .A1(n1592), .B0(n1578), .B1(n4848), .C0(n1564), 
        .C1(n4847), .Y(n3777) );
  INVX1 U4408 ( .A(prev_key0_reg[7]), .Y(n4847) );
  INVX1 U4409 ( .A(sboxw[7]), .Y(n4848) );
  OAI222XL U4410 ( .A0(n5789), .A1(n1591), .B0(n1577), .B1(n4881), .C0(n1557), 
        .C1(n4880), .Y(n3776) );
  INVX1 U4411 ( .A(prev_key0_reg[8]), .Y(n4880) );
  INVX1 U4412 ( .A(sboxw[8]), .Y(n4881) );
  OAI222XL U4413 ( .A0(n5773), .A1(n1594), .B0(n1578), .B1(n4914), .C0(n1563), 
        .C1(n4913), .Y(n3775) );
  INVX1 U4414 ( .A(prev_key0_reg[9]), .Y(n4913) );
  INVX1 U4415 ( .A(sboxw[9]), .Y(n4914) );
  OAI222XL U4416 ( .A0(n5805), .A1(n1593), .B0(n1577), .B1(n4947), .C0(n1564), 
        .C1(n4946), .Y(n3774) );
  INVX1 U4417 ( .A(prev_key0_reg[10]), .Y(n4946) );
  INVX1 U4418 ( .A(sboxw[10]), .Y(n4947) );
  OAI222XL U4419 ( .A0(n5821), .A1(n1590), .B0(n1567), .B1(n4980), .C0(n1557), 
        .C1(n4979), .Y(n3773) );
  INVX1 U4420 ( .A(prev_key0_reg[11]), .Y(n4979) );
  INVX1 U4421 ( .A(sboxw[11]), .Y(n4980) );
  OAI222XL U4422 ( .A0(n5837), .A1(n1582), .B0(n1567), .B1(n5013), .C0(n1562), 
        .C1(n5012), .Y(n3772) );
  INVX1 U4423 ( .A(prev_key0_reg[12]), .Y(n5012) );
  INVX1 U4424 ( .A(sboxw[12]), .Y(n5013) );
  OAI222XL U4425 ( .A0(n5853), .A1(n1582), .B0(n1580), .B1(n5046), .C0(n1564), 
        .C1(n5045), .Y(n3771) );
  INVX1 U4426 ( .A(prev_key0_reg[13]), .Y(n5045) );
  INVX1 U4427 ( .A(sboxw[13]), .Y(n5046) );
  OAI222XL U4428 ( .A0(n5869), .A1(n1582), .B0(n1580), .B1(n5078), .C0(n1566), 
        .C1(n5077), .Y(n3770) );
  INVX1 U4429 ( .A(prev_key0_reg[14]), .Y(n5077) );
  INVX1 U4430 ( .A(sboxw[14]), .Y(n5078) );
  OAI222XL U4431 ( .A0(n5885), .A1(n1583), .B0(n1580), .B1(n5111), .C0(n1564), 
        .C1(n5110), .Y(n3769) );
  INVX1 U4432 ( .A(prev_key0_reg[15]), .Y(n5110) );
  INVX1 U4433 ( .A(sboxw[15]), .Y(n5111) );
  OAI222XL U4434 ( .A0(n5791), .A1(n1583), .B0(n1569), .B1(n5144), .C0(n1566), 
        .C1(n5143), .Y(n3768) );
  INVX1 U4435 ( .A(prev_key0_reg[16]), .Y(n5143) );
  INVX1 U4436 ( .A(sboxw[16]), .Y(n5144) );
  OAI222XL U4437 ( .A0(n5779), .A1(n1584), .B0(n1569), .B1(n5177), .C0(n1565), 
        .C1(n5176), .Y(n3767) );
  INVX1 U4438 ( .A(prev_key0_reg[17]), .Y(n5176) );
  INVX1 U4439 ( .A(sboxw[17]), .Y(n5177) );
  OAI222XL U4440 ( .A0(n5807), .A1(n1584), .B0(n1569), .B1(n5210), .C0(n1556), 
        .C1(n5209), .Y(n3766) );
  INVX1 U4441 ( .A(prev_key0_reg[18]), .Y(n5209) );
  INVX1 U4442 ( .A(sboxw[18]), .Y(n5210) );
  OAI222XL U4443 ( .A0(n5823), .A1(n1584), .B0(n1576), .B1(n5243), .C0(n1556), 
        .C1(n5242), .Y(n3765) );
  INVX1 U4444 ( .A(prev_key0_reg[19]), .Y(n5242) );
  INVX1 U4445 ( .A(sboxw[19]), .Y(n5243) );
  OAI222XL U4446 ( .A0(n5839), .A1(n1585), .B0(n1576), .B1(n5276), .C0(n1556), 
        .C1(n5275), .Y(n3764) );
  INVX1 U4447 ( .A(prev_key0_reg[20]), .Y(n5275) );
  INVX1 U4448 ( .A(sboxw[20]), .Y(n5276) );
  OAI222XL U4449 ( .A0(n5855), .A1(n1585), .B0(n1576), .B1(n5309), .C0(n1562), 
        .C1(n5308), .Y(n3763) );
  INVX1 U4450 ( .A(prev_key0_reg[21]), .Y(n5308) );
  INVX1 U4451 ( .A(sboxw[21]), .Y(n5309) );
  OAI222XL U4452 ( .A0(n5871), .A1(n1586), .B0(n1575), .B1(n5341), .C0(n1563), 
        .C1(n5340), .Y(n3762) );
  INVX1 U4453 ( .A(prev_key0_reg[22]), .Y(n5340) );
  INVX1 U4454 ( .A(sboxw[22]), .Y(n5341) );
  OAI222XL U4455 ( .A0(n5887), .A1(n1586), .B0(n1569), .B1(n5374), .C0(n1562), 
        .C1(n5373), .Y(n3761) );
  INVX1 U4456 ( .A(prev_key0_reg[23]), .Y(n5373) );
  INVX1 U4457 ( .A(sboxw[23]), .Y(n5374) );
  OAI222XL U4458 ( .A0(n5792), .A1(n1581), .B0(n1568), .B1(n4623), .C0(n1559), 
        .C1(n4622), .Y(n3752) );
  INVX1 U4459 ( .A(prev_key0_reg[32]), .Y(n4622) );
  INVX1 U4460 ( .A(prev_key1_reg[32]), .Y(n4623) );
  OAI222XL U4461 ( .A0(n5775), .A1(n1581), .B0(n1577), .B1(n4655), .C0(n1558), 
        .C1(n4654), .Y(n3751) );
  INVX1 U4462 ( .A(prev_key0_reg[33]), .Y(n4654) );
  INVX1 U4463 ( .A(prev_key1_reg[33]), .Y(n4655) );
  OAI222XL U4464 ( .A0(n5808), .A1(n1594), .B0(n1579), .B1(n4687), .C0(n1559), 
        .C1(n4686), .Y(n3750) );
  INVX1 U4465 ( .A(prev_key0_reg[34]), .Y(n4686) );
  INVX1 U4466 ( .A(prev_key1_reg[34]), .Y(n4687) );
  OAI222XL U4467 ( .A0(n5824), .A1(n1593), .B0(n1568), .B1(n4719), .C0(n1558), 
        .C1(n4718), .Y(n3749) );
  INVX1 U4468 ( .A(prev_key0_reg[35]), .Y(n4718) );
  INVX1 U4469 ( .A(prev_key1_reg[35]), .Y(n4719) );
  OAI222XL U4470 ( .A0(n5840), .A1(n1590), .B0(n1568), .B1(n4751), .C0(n1558), 
        .C1(n4750), .Y(n3748) );
  INVX1 U4471 ( .A(prev_key0_reg[36]), .Y(n4750) );
  INVX1 U4472 ( .A(prev_key1_reg[36]), .Y(n4751) );
  OAI222XL U4473 ( .A0(n5856), .A1(n1593), .B0(n5661), .B1(n4783), .C0(n1558), 
        .C1(n4782), .Y(n3747) );
  INVX1 U4474 ( .A(prev_key0_reg[37]), .Y(n4782) );
  INVX1 U4475 ( .A(prev_key1_reg[37]), .Y(n4783) );
  OAI222XL U4476 ( .A0(n5872), .A1(n1590), .B0(n1579), .B1(n4814), .C0(n1557), 
        .C1(n4813), .Y(n3746) );
  INVX1 U4477 ( .A(prev_key0_reg[38]), .Y(n4813) );
  INVX1 U4478 ( .A(prev_key1_reg[38]), .Y(n4814) );
  OAI222XL U4479 ( .A0(n5888), .A1(n5663), .B0(n1568), .B1(n4846), .C0(n1558), 
        .C1(n4845), .Y(n3745) );
  INVX1 U4480 ( .A(prev_key0_reg[39]), .Y(n4845) );
  INVX1 U4481 ( .A(prev_key1_reg[39]), .Y(n4846) );
  OAI222XL U4482 ( .A0(n5787), .A1(n5663), .B0(n1568), .B1(n4879), .C0(n1565), 
        .C1(n4878), .Y(n3744) );
  INVX1 U4483 ( .A(prev_key0_reg[40]), .Y(n4878) );
  INVX1 U4484 ( .A(prev_key1_reg[40]), .Y(n4879) );
  OAI222XL U4485 ( .A0(n5767), .A1(n1592), .B0(n5661), .B1(n4912), .C0(n1564), 
        .C1(n4911), .Y(n3743) );
  INVX1 U4486 ( .A(prev_key0_reg[41]), .Y(n4911) );
  INVX1 U4487 ( .A(prev_key1_reg[41]), .Y(n4912) );
  OAI222XL U4488 ( .A0(n5803), .A1(n1592), .B0(n1578), .B1(n4945), .C0(n1561), 
        .C1(n4944), .Y(n3742) );
  INVX1 U4489 ( .A(prev_key0_reg[42]), .Y(n4944) );
  INVX1 U4490 ( .A(prev_key1_reg[42]), .Y(n4945) );
  OAI222XL U4491 ( .A0(n5819), .A1(n1591), .B0(n1577), .B1(n4978), .C0(n1557), 
        .C1(n4977), .Y(n3741) );
  INVX1 U4492 ( .A(prev_key0_reg[43]), .Y(n4977) );
  INVX1 U4493 ( .A(prev_key1_reg[43]), .Y(n4978) );
  OAI222XL U4494 ( .A0(n5835), .A1(n1582), .B0(n1567), .B1(n5011), .C0(n1557), 
        .C1(n5010), .Y(n3740) );
  INVX1 U4495 ( .A(prev_key0_reg[44]), .Y(n5010) );
  INVX1 U4496 ( .A(prev_key1_reg[44]), .Y(n5011) );
  OAI222XL U4497 ( .A0(n5851), .A1(n1582), .B0(n1580), .B1(n5044), .C0(n1565), 
        .C1(n5043), .Y(n3739) );
  INVX1 U4498 ( .A(prev_key0_reg[45]), .Y(n5043) );
  INVX1 U4499 ( .A(prev_key1_reg[45]), .Y(n5044) );
  OAI222XL U4500 ( .A0(n5867), .A1(n1582), .B0(n1580), .B1(n5076), .C0(n1566), 
        .C1(n5075), .Y(n3738) );
  INVX1 U4501 ( .A(prev_key0_reg[46]), .Y(n5075) );
  INVX1 U4502 ( .A(prev_key1_reg[46]), .Y(n5076) );
  OAI222XL U4503 ( .A0(n5883), .A1(n1583), .B0(n1580), .B1(n5109), .C0(n1566), 
        .C1(n5108), .Y(n3737) );
  INVX1 U4504 ( .A(prev_key0_reg[47]), .Y(n5108) );
  INVX1 U4505 ( .A(prev_key1_reg[47]), .Y(n5109) );
  OAI222XL U4506 ( .A0(n5793), .A1(n1583), .B0(n1569), .B1(n5142), .C0(n1565), 
        .C1(n5141), .Y(n3736) );
  INVX1 U4507 ( .A(prev_key0_reg[48]), .Y(n5141) );
  INVX1 U4508 ( .A(prev_key1_reg[48]), .Y(n5142) );
  OAI222XL U4509 ( .A0(n5777), .A1(n1584), .B0(n1569), .B1(n5175), .C0(n1564), 
        .C1(n5174), .Y(n3735) );
  INVX1 U4510 ( .A(prev_key0_reg[49]), .Y(n5174) );
  INVX1 U4511 ( .A(prev_key1_reg[49]), .Y(n5175) );
  OAI222XL U4512 ( .A0(n5809), .A1(n1584), .B0(n1569), .B1(n5208), .C0(n1556), 
        .C1(n5207), .Y(n3734) );
  INVX1 U4513 ( .A(prev_key0_reg[50]), .Y(n5207) );
  INVX1 U4514 ( .A(prev_key1_reg[50]), .Y(n5208) );
  OAI222XL U4515 ( .A0(n5825), .A1(n1584), .B0(n1576), .B1(n5241), .C0(n1556), 
        .C1(n5240), .Y(n3733) );
  INVX1 U4516 ( .A(prev_key0_reg[51]), .Y(n5240) );
  INVX1 U4517 ( .A(prev_key1_reg[51]), .Y(n5241) );
  OAI222XL U4518 ( .A0(n5841), .A1(n1585), .B0(n1576), .B1(n5274), .C0(n1556), 
        .C1(n5273), .Y(n3732) );
  INVX1 U4519 ( .A(prev_key0_reg[52]), .Y(n5273) );
  INVX1 U4520 ( .A(prev_key1_reg[52]), .Y(n5274) );
  OAI222XL U4521 ( .A0(n5857), .A1(n1585), .B0(n1576), .B1(n5307), .C0(n1562), 
        .C1(n5306), .Y(n3731) );
  INVX1 U4522 ( .A(prev_key0_reg[53]), .Y(n5306) );
  INVX1 U4523 ( .A(prev_key1_reg[53]), .Y(n5307) );
  OAI222XL U4524 ( .A0(n5873), .A1(n1586), .B0(n1575), .B1(n5339), .C0(n1563), 
        .C1(n5338), .Y(n3730) );
  INVX1 U4525 ( .A(prev_key0_reg[54]), .Y(n5338) );
  INVX1 U4526 ( .A(prev_key1_reg[54]), .Y(n5339) );
  OAI222XL U4527 ( .A0(n5889), .A1(n1586), .B0(n1575), .B1(n5372), .C0(n1), 
        .C1(n5371), .Y(n3729) );
  INVX1 U4528 ( .A(prev_key0_reg[55]), .Y(n5371) );
  INVX1 U4529 ( .A(prev_key1_reg[55]), .Y(n5372) );
  OAI222XL U4530 ( .A0(n5796), .A1(n1581), .B0(n1572), .B1(n4590), .C0(n1553), 
        .C1(n4609), .Y(n3688) );
  INVX1 U4531 ( .A(prev_key1_reg[96]), .Y(n4590) );
  OAI222XL U4532 ( .A0(n5774), .A1(n1581), .B0(n1567), .B1(n4634), .C0(n1559), 
        .C1(n4640), .Y(n3687) );
  INVX1 U4533 ( .A(prev_key1_reg[97]), .Y(n4634) );
  OAI222XL U4534 ( .A0(n5812), .A1(n1581), .B0(n1578), .B1(n4666), .C0(n1559), 
        .C1(n4672), .Y(n3913) );
  INVX1 U4535 ( .A(prev_key1_reg[98]), .Y(n4666) );
  OAI222XL U4536 ( .A0(n5828), .A1(n1592), .B0(n5661), .B1(n4698), .C0(n1558), 
        .C1(n4704), .Y(n3686) );
  INVX1 U4537 ( .A(prev_key1_reg[99]), .Y(n4698) );
  OAI222XL U4538 ( .A0(n5844), .A1(n1591), .B0(n5661), .B1(n4730), .C0(n1558), 
        .C1(n4736), .Y(n3685) );
  INVX1 U4539 ( .A(prev_key1_reg[100]), .Y(n4730) );
  OAI222XL U4540 ( .A0(n5860), .A1(n1592), .B0(n5661), .B1(n4762), .C0(n1558), 
        .C1(n4768), .Y(n3684) );
  INVX1 U4541 ( .A(prev_key1_reg[101]), .Y(n4762) );
  OAI222XL U4542 ( .A0(n5892), .A1(n1591), .B0(n5661), .B1(n4825), .C0(n1558), 
        .C1(n4831), .Y(n3682) );
  INVX1 U4543 ( .A(prev_key1_reg[103]), .Y(n4825) );
  OAI222XL U4544 ( .A0(n5783), .A1(n1591), .B0(n1579), .B1(n4857), .C0(n1566), 
        .C1(n4864), .Y(n3681) );
  INVX1 U4545 ( .A(prev_key1_reg[104]), .Y(n4857) );
  OAI222XL U4546 ( .A0(n5766), .A1(n1594), .B0(n1578), .B1(n4890), .C0(n1557), 
        .C1(n4897), .Y(n3680) );
  INVX1 U4547 ( .A(prev_key1_reg[105]), .Y(n4890) );
  OAI222XL U4548 ( .A0(n5799), .A1(n1594), .B0(n1578), .B1(n4923), .C0(n1564), 
        .C1(n4930), .Y(n3679) );
  INVX1 U4549 ( .A(prev_key1_reg[106]), .Y(n4923) );
  OAI222XL U4550 ( .A0(n5815), .A1(n5663), .B0(n1577), .B1(n4956), .C0(n1557), 
        .C1(n4963), .Y(n3678) );
  INVX1 U4551 ( .A(prev_key1_reg[107]), .Y(n4956) );
  OAI222XL U4552 ( .A0(n5831), .A1(n1590), .B0(n1567), .B1(n4989), .C0(n1564), 
        .C1(n4996), .Y(n3677) );
  INVX1 U4553 ( .A(prev_key1_reg[108]), .Y(n4989) );
  OAI222XL U4554 ( .A0(n5847), .A1(n1582), .B0(n1580), .B1(n5022), .C0(n1562), 
        .C1(n5029), .Y(n3676) );
  INVX1 U4555 ( .A(prev_key1_reg[109]), .Y(n5022) );
  OAI222XL U4556 ( .A0(n5863), .A1(n1582), .B0(n1568), .B1(n5055), .C0(n1561), 
        .C1(n5062), .Y(n3675) );
  INVX1 U4557 ( .A(prev_key1_reg[110]), .Y(n5055) );
  OAI222XL U4558 ( .A0(n5879), .A1(n1583), .B0(n1580), .B1(n5087), .C0(n1563), 
        .C1(n5094), .Y(n3674) );
  INVX1 U4559 ( .A(prev_key1_reg[111]), .Y(n5087) );
  OAI222XL U4560 ( .A0(n5797), .A1(n1583), .B0(n1567), .B1(n5120), .C0(n1566), 
        .C1(n5127), .Y(n3673) );
  INVX1 U4561 ( .A(prev_key1_reg[112]), .Y(n5120) );
  OAI222XL U4562 ( .A0(n5776), .A1(n1583), .B0(n1569), .B1(n5153), .C0(n1565), 
        .C1(n5160), .Y(n3672) );
  INVX1 U4563 ( .A(prev_key1_reg[113]), .Y(n5153) );
  OAI222XL U4564 ( .A0(n5813), .A1(n1584), .B0(n1580), .B1(n5186), .C0(n1556), 
        .C1(n5193), .Y(n3671) );
  INVX1 U4565 ( .A(prev_key1_reg[114]), .Y(n5186) );
  OAI222XL U4566 ( .A0(n5829), .A1(n1584), .B0(n1576), .B1(n5219), .C0(n1556), 
        .C1(n5226), .Y(n3670) );
  INVX1 U4567 ( .A(prev_key1_reg[115]), .Y(n5219) );
  OAI222XL U4568 ( .A0(n5845), .A1(n1585), .B0(n1576), .B1(n5252), .C0(n1556), 
        .C1(n5259), .Y(n3669) );
  INVX1 U4569 ( .A(prev_key1_reg[116]), .Y(n5252) );
  OAI222XL U4570 ( .A0(n5861), .A1(n1585), .B0(n1576), .B1(n5285), .C0(n1556), 
        .C1(n5292), .Y(n3668) );
  INVX1 U4571 ( .A(prev_key1_reg[117]), .Y(n5285) );
  OAI222XL U4572 ( .A0(n5877), .A1(n1585), .B0(n1576), .B1(n5318), .C0(n1), 
        .C1(n5325), .Y(n3667) );
  INVX1 U4573 ( .A(prev_key1_reg[118]), .Y(n5318) );
  OAI222XL U4574 ( .A0(n5893), .A1(n1586), .B0(n1575), .B1(n5350), .C0(n1), 
        .C1(n5357), .Y(n3666) );
  INVX1 U4575 ( .A(prev_key1_reg[119]), .Y(n5350) );
  OAI222XL U4576 ( .A0(n5794), .A1(n1581), .B0(n194), .B1(n1561), .C0(n1570), 
        .C1(n4615), .Y(n3720) );
  INVX1 U4577 ( .A(prev_key1_reg[64]), .Y(n4615) );
  OAI222XL U4578 ( .A0(n5780), .A1(n1581), .B0(n193), .B1(n1561), .C0(n1570), 
        .C1(n4646), .Y(n3719) );
  INVX1 U4579 ( .A(prev_key1_reg[65]), .Y(n4646) );
  OAI222XL U4580 ( .A0(n5810), .A1(n1581), .B0(n192), .B1(n1561), .C0(n1570), 
        .C1(n4678), .Y(n3718) );
  INVX1 U4581 ( .A(prev_key1_reg[66]), .Y(n4678) );
  OAI222XL U4582 ( .A0(n5826), .A1(n1593), .B0(n191), .B1(n1561), .C0(n1570), 
        .C1(n4710), .Y(n3717) );
  INVX1 U4583 ( .A(prev_key1_reg[67]), .Y(n4710) );
  OAI222XL U4584 ( .A0(n5842), .A1(n1593), .B0(n190), .B1(n1561), .C0(n1570), 
        .C1(n4742), .Y(n3716) );
  INVX1 U4585 ( .A(prev_key1_reg[68]), .Y(n4742) );
  OAI222XL U4586 ( .A0(n5858), .A1(n1590), .B0(n189), .B1(n1561), .C0(n1570), 
        .C1(n4774), .Y(n3715) );
  INVX1 U4587 ( .A(prev_key1_reg[69]), .Y(n4774) );
  OAI222XL U4588 ( .A0(n5874), .A1(n1592), .B0(n188), .B1(n1561), .C0(n1571), 
        .C1(n4805), .Y(n3714) );
  INVX1 U4589 ( .A(prev_key1_reg[70]), .Y(n4805) );
  OAI222XL U4590 ( .A0(n5890), .A1(n1593), .B0(n187), .B1(n1560), .C0(n1571), 
        .C1(n4837), .Y(n3713) );
  INVX1 U4591 ( .A(prev_key1_reg[71]), .Y(n4837) );
  OAI222XL U4592 ( .A0(n5785), .A1(n1590), .B0(n186), .B1(n1560), .C0(n1571), 
        .C1(n4870), .Y(n3712) );
  INVX1 U4593 ( .A(prev_key1_reg[72]), .Y(n4870) );
  OAI222XL U4594 ( .A0(n5772), .A1(n1593), .B0(n185), .B1(n1559), .C0(n1571), 
        .C1(n4903), .Y(n3711) );
  INVX1 U4595 ( .A(prev_key1_reg[73]), .Y(n4903) );
  OAI222XL U4596 ( .A0(n5801), .A1(n1589), .B0(n184), .B1(n1559), .C0(n1571), 
        .C1(n4936), .Y(n3710) );
  INVX1 U4597 ( .A(prev_key1_reg[74]), .Y(n4936) );
  OAI222XL U4598 ( .A0(n5817), .A1(n1589), .B0(n183), .B1(n1560), .C0(n1571), 
        .C1(n4969), .Y(n3709) );
  INVX1 U4599 ( .A(prev_key1_reg[75]), .Y(n4969) );
  OAI222XL U4600 ( .A0(n5833), .A1(n1593), .B0(n182), .B1(n1559), .C0(n1571), 
        .C1(n5002), .Y(n3708) );
  INVX1 U4601 ( .A(prev_key1_reg[76]), .Y(n5002) );
  OAI222XL U4602 ( .A0(n5849), .A1(n1582), .B0(n181), .B1(n1559), .C0(n1571), 
        .C1(n5035), .Y(n3707) );
  INVX1 U4603 ( .A(prev_key1_reg[77]), .Y(n5035) );
  OAI222XL U4604 ( .A0(n5865), .A1(n1582), .B0(n180), .B1(n1559), .C0(n1571), 
        .C1(n5067), .Y(n3706) );
  INVX1 U4605 ( .A(prev_key1_reg[78]), .Y(n5067) );
  OAI222XL U4606 ( .A0(n5881), .A1(n1583), .B0(n179), .B1(n1559), .C0(n1572), 
        .C1(n5100), .Y(n3705) );
  INVX1 U4607 ( .A(prev_key1_reg[79]), .Y(n5100) );
  OAI222XL U4608 ( .A0(n5795), .A1(n1583), .B0(n178), .B1(n1560), .C0(n1572), 
        .C1(n5133), .Y(n3704) );
  INVX1 U4609 ( .A(prev_key1_reg[80]), .Y(n5133) );
  OAI222XL U4610 ( .A0(n5778), .A1(n1583), .B0(n177), .B1(n1560), .C0(n1572), 
        .C1(n5166), .Y(n3703) );
  INVX1 U4611 ( .A(prev_key1_reg[81]), .Y(n5166) );
  OAI222XL U4612 ( .A0(n5811), .A1(n1584), .B0(n176), .B1(n1560), .C0(n1570), 
        .C1(n5199), .Y(n3702) );
  INVX1 U4613 ( .A(prev_key1_reg[82]), .Y(n5199) );
  OAI222XL U4614 ( .A0(n5827), .A1(n1584), .B0(n175), .B1(n1561), .C0(n1572), 
        .C1(n5232), .Y(n3701) );
  INVX1 U4615 ( .A(prev_key1_reg[83]), .Y(n5232) );
  OAI222XL U4616 ( .A0(n5843), .A1(n1585), .B0(n174), .B1(n1560), .C0(n1570), 
        .C1(n5265), .Y(n3700) );
  INVX1 U4617 ( .A(prev_key1_reg[84]), .Y(n5265) );
  OAI222XL U4618 ( .A0(n5859), .A1(n1585), .B0(n173), .B1(n1560), .C0(n1570), 
        .C1(n5298), .Y(n3699) );
  INVX1 U4619 ( .A(prev_key1_reg[85]), .Y(n5298) );
  OAI222XL U4620 ( .A0(n5875), .A1(n1585), .B0(n172), .B1(n1560), .C0(n1571), 
        .C1(n5331), .Y(n3698) );
  INVX1 U4621 ( .A(prev_key1_reg[86]), .Y(n5331) );
  OAI222XL U4622 ( .A0(n5891), .A1(n1586), .B0(n171), .B1(n1560), .C0(n1570), 
        .C1(n5363), .Y(n3697) );
  INVX1 U4623 ( .A(prev_key1_reg[87]), .Y(n5363) );
  OAI222XL U4624 ( .A0(n5876), .A1(n1594), .B0(n5661), .B1(n4794), .C0(n1558), 
        .C1(n4799), .Y(n3683) );
  INVX1 U4625 ( .A(prev_key1_reg[102]), .Y(n4794) );
  OAI221XL U4626 ( .A0(n1668), .A1(n4995), .B0(n4994), .B1(n1657), .C0(n4993), 
        .Y(n3804) );
  INVX1 U4627 ( .A(key[108]), .Y(n4995) );
  AOI221XL U4628 ( .A0(n1642), .A1(n823), .B0(n1632), .B1(key[236]), .C0(n4992), .Y(n4993) );
  MXI4X1 U4629 ( .A(n246), .B(n247), .C(n248), .D(n249), .S0(n1271), .S1(n1286), .Y(round_key[29]) );
  MXI4X1 U4630 ( .A(\key_mem[4][29] ), .B(\key_mem[5][29] ), .C(
        \key_mem[6][29] ), .D(\key_mem[7][29] ), .S0(n1359), .S1(n1332), .Y(
        n248) );
  MXI3X1 U4631 ( .A(\key_mem[12][29] ), .B(\key_mem[13][29] ), .C(n245), .S0(
        n1372), .S1(n1339), .Y(n249) );
  MXI4X1 U4632 ( .A(\key_mem[0][29] ), .B(\key_mem[1][29] ), .C(
        \key_mem[2][29] ), .D(\key_mem[3][29] ), .S0(n1417), .S1(n1333), .Y(
        n246) );
  MXI4X1 U4633 ( .A(n241), .B(n242), .C(n243), .D(n244), .S0(n1271), .S1(n1286), .Y(round_key[28]) );
  MXI4X1 U4634 ( .A(\key_mem[4][28] ), .B(\key_mem[5][28] ), .C(
        \key_mem[6][28] ), .D(\key_mem[7][28] ), .S0(n1352), .S1(n1331), .Y(
        n243) );
  MXI3X1 U4635 ( .A(\key_mem[12][28] ), .B(\key_mem[13][28] ), .C(n240), .S0(
        n1372), .S1(n1339), .Y(n244) );
  MXI4X1 U4636 ( .A(\key_mem[0][28] ), .B(\key_mem[1][28] ), .C(
        \key_mem[2][28] ), .D(\key_mem[3][28] ), .S0(N31), .S1(n1333), .Y(n241) );
  MXI4X1 U4637 ( .A(n236), .B(n237), .C(n238), .D(n239), .S0(n1270), .S1(n1285), .Y(round_key[27]) );
  MXI4X1 U4638 ( .A(\key_mem[4][27] ), .B(\key_mem[5][27] ), .C(
        \key_mem[6][27] ), .D(\key_mem[7][27] ), .S0(n1415), .S1(n1333), .Y(
        n238) );
  MXI3X1 U4639 ( .A(\key_mem[12][27] ), .B(\key_mem[13][27] ), .C(n235), .S0(
        n1371), .S1(n1339), .Y(n239) );
  MXI4X1 U4640 ( .A(\key_mem[0][27] ), .B(\key_mem[1][27] ), .C(
        \key_mem[2][27] ), .D(\key_mem[3][27] ), .S0(n1368), .S1(n1333), .Y(
        n236) );
  MXI4X1 U4641 ( .A(n231), .B(n232), .C(n233), .D(n234), .S0(n1270), .S1(n1285), .Y(round_key[26]) );
  MXI4X1 U4642 ( .A(\key_mem[4][26] ), .B(\key_mem[5][26] ), .C(
        \key_mem[6][26] ), .D(\key_mem[7][26] ), .S0(n1410), .S1(n1334), .Y(
        n233) );
  MXI3X1 U4643 ( .A(\key_mem[12][26] ), .B(\key_mem[13][26] ), .C(n230), .S0(
        n1371), .S1(n1339), .Y(n234) );
  MXI4X1 U4644 ( .A(\key_mem[0][26] ), .B(\key_mem[1][26] ), .C(
        \key_mem[2][26] ), .D(\key_mem[3][26] ), .S0(n1410), .S1(n1332), .Y(
        n231) );
  MXI4X1 U4645 ( .A(n395), .B(n396), .C(n397), .D(n398), .S0(n1273), .S1(n1288), .Y(round_key[56]) );
  MXI4X1 U4646 ( .A(\key_mem[4][56] ), .B(\key_mem[5][56] ), .C(
        \key_mem[6][56] ), .D(\key_mem[7][56] ), .S0(n1381), .S1(n1312), .Y(
        n397) );
  MXI3X1 U4647 ( .A(\key_mem[12][56] ), .B(\key_mem[13][56] ), .C(n394), .S0(
        n1377), .S1(n1342), .Y(n398) );
  MXI4X1 U4648 ( .A(\key_mem[0][56] ), .B(\key_mem[1][56] ), .C(
        \key_mem[2][56] ), .D(\key_mem[3][56] ), .S0(n1382), .S1(n1312), .Y(
        n395) );
  MXI4X1 U4649 ( .A(n420), .B(n421), .C(n422), .D(n423), .S0(n1269), .S1(n1282), .Y(round_key[61]) );
  MXI4X1 U4650 ( .A(\key_mem[4][61] ), .B(\key_mem[5][61] ), .C(
        \key_mem[6][61] ), .D(\key_mem[7][61] ), .S0(n1385), .S1(n1314), .Y(
        n422) );
  MXI3X1 U4651 ( .A(\key_mem[12][61] ), .B(\key_mem[13][61] ), .C(n419), .S0(
        n1380), .S1(n1342), .Y(n423) );
  MXI4X1 U4652 ( .A(\key_mem[0][61] ), .B(\key_mem[1][61] ), .C(
        \key_mem[2][61] ), .D(\key_mem[3][61] ), .S0(n1385), .S1(n1314), .Y(
        n420) );
  MXI4X1 U4653 ( .A(n415), .B(n416), .C(n417), .D(n418), .S0(n1267), .S1(n1290), .Y(round_key[60]) );
  MXI4X1 U4654 ( .A(\key_mem[4][60] ), .B(\key_mem[5][60] ), .C(
        \key_mem[6][60] ), .D(\key_mem[7][60] ), .S0(n1384), .S1(n1313), .Y(
        n417) );
  MXI3X1 U4655 ( .A(\key_mem[12][60] ), .B(\key_mem[13][60] ), .C(n414), .S0(
        n1380), .S1(n1342), .Y(n418) );
  MXI4X1 U4656 ( .A(\key_mem[0][60] ), .B(\key_mem[1][60] ), .C(
        \key_mem[2][60] ), .D(\key_mem[3][60] ), .S0(n1384), .S1(n1314), .Y(
        n415) );
  MXI4X1 U4657 ( .A(n400), .B(n401), .C(n402), .D(n403), .S0(n1273), .S1(n1288), .Y(round_key[57]) );
  MXI4X1 U4658 ( .A(\key_mem[4][57] ), .B(\key_mem[5][57] ), .C(
        \key_mem[6][57] ), .D(\key_mem[7][57] ), .S0(n1382), .S1(n1312), .Y(
        n402) );
  MXI3X1 U4659 ( .A(\key_mem[12][57] ), .B(\key_mem[13][57] ), .C(n399), .S0(
        n1379), .S1(n1342), .Y(n403) );
  MXI4X1 U4660 ( .A(\key_mem[0][57] ), .B(\key_mem[1][57] ), .C(
        \key_mem[2][57] ), .D(\key_mem[3][57] ), .S0(n1382), .S1(n1312), .Y(
        n400) );
  MXI4X1 U4661 ( .A(n221), .B(n222), .C(n223), .D(n224), .S0(n1270), .S1(n1285), .Y(round_key[24]) );
  MXI3X1 U4662 ( .A(\key_mem[12][24] ), .B(\key_mem[13][24] ), .C(n220), .S0(
        n1370), .S1(n1339), .Y(n224) );
  MXI4X1 U4663 ( .A(\key_mem[4][24] ), .B(\key_mem[5][24] ), .C(
        \key_mem[6][24] ), .D(\key_mem[7][24] ), .S0(n1410), .S1(n1296), .Y(
        n223) );
  MXI4X1 U4664 ( .A(\key_mem[0][24] ), .B(\key_mem[1][24] ), .C(
        \key_mem[2][24] ), .D(\key_mem[3][24] ), .S0(n1410), .S1(n1306), .Y(
        n221) );
  MXI4X1 U4665 ( .A(n256), .B(n257), .C(n258), .D(n259), .S0(n1271), .S1(n1286), .Y(round_key[31]) );
  MXI4X1 U4666 ( .A(\key_mem[4][31] ), .B(\key_mem[5][31] ), .C(
        \key_mem[6][31] ), .D(\key_mem[7][31] ), .S0(n1356), .S1(n1333), .Y(
        n258) );
  MXI3X1 U4667 ( .A(\key_mem[12][31] ), .B(\key_mem[13][31] ), .C(n255), .S0(
        n1373), .S1(n1339), .Y(n259) );
  MXI4X1 U4668 ( .A(\key_mem[0][31] ), .B(\key_mem[1][31] ), .C(
        \key_mem[2][31] ), .D(\key_mem[3][31] ), .S0(n1351), .S1(n1332), .Y(
        n256) );
  MXI4X1 U4669 ( .A(n251), .B(n252), .C(n253), .D(n254), .S0(n1271), .S1(n1286), .Y(round_key[30]) );
  MXI4X1 U4670 ( .A(\key_mem[4][30] ), .B(\key_mem[5][30] ), .C(
        \key_mem[6][30] ), .D(\key_mem[7][30] ), .S0(n1361), .S1(n1331), .Y(
        n253) );
  MXI3X1 U4671 ( .A(\key_mem[12][30] ), .B(\key_mem[13][30] ), .C(n250), .S0(
        n1373), .S1(n1339), .Y(n254) );
  MXI4X1 U4672 ( .A(\key_mem[0][30] ), .B(\key_mem[1][30] ), .C(
        \key_mem[2][30] ), .D(\key_mem[3][30] ), .S0(n1365), .S1(n1332), .Y(
        n251) );
  MXI4X1 U4673 ( .A(n1256), .B(n1257), .C(n1258), .D(n1259), .S0(n1276), .S1(
        n1289), .Y(round_key[126]) );
  MXI4X1 U4674 ( .A(\key_mem[4][126] ), .B(\key_mem[5][126] ), .C(
        \key_mem[6][126] ), .D(\key_mem[7][126] ), .S0(n1388), .S1(n1302), .Y(
        n1258) );
  MXI3X1 U4675 ( .A(\key_mem[12][126] ), .B(\key_mem[13][126] ), .C(n1255), 
        .S0(n1377), .S1(n1335), .Y(n1259) );
  MXI4X1 U4676 ( .A(\key_mem[0][126] ), .B(\key_mem[1][126] ), .C(
        \key_mem[2][126] ), .D(\key_mem[3][126] ), .S0(n1388), .S1(n1298), .Y(
        n1256) );
  MXI4X1 U4677 ( .A(n1248), .B(n1251), .C(n1252), .D(n1253), .S0(n1276), .S1(
        n1289), .Y(round_key[125]) );
  MXI4X1 U4678 ( .A(\key_mem[4][125] ), .B(\key_mem[5][125] ), .C(
        \key_mem[6][125] ), .D(\key_mem[7][125] ), .S0(n1389), .S1(n1305), .Y(
        n1252) );
  MXI3X1 U4679 ( .A(\key_mem[12][125] ), .B(\key_mem[13][125] ), .C(n1247), 
        .S0(n1377), .S1(n1335), .Y(n1253) );
  MXI4X1 U4680 ( .A(\key_mem[0][125] ), .B(\key_mem[1][125] ), .C(
        \key_mem[2][125] ), .D(\key_mem[3][125] ), .S0(n1389), .S1(n1305), .Y(
        n1248) );
  MXI4X1 U4681 ( .A(n1208), .B(n1211), .C(n1212), .D(n1215), .S0(n1276), .S1(
        n1289), .Y(round_key[121]) );
  MXI4X1 U4682 ( .A(\key_mem[4][121] ), .B(\key_mem[5][121] ), .C(
        \key_mem[6][121] ), .D(\key_mem[7][121] ), .S0(n1390), .S1(n1300), .Y(
        n1212) );
  MXI3X1 U4683 ( .A(\key_mem[12][121] ), .B(\key_mem[13][121] ), .C(n1207), 
        .S0(n1380), .S1(n1336), .Y(n1215) );
  MXI4X1 U4684 ( .A(\key_mem[0][121] ), .B(\key_mem[1][121] ), .C(
        \key_mem[2][121] ), .D(\key_mem[3][121] ), .S0(n1390), .S1(n1294), .Y(
        n1208) );
  MXI4X1 U4685 ( .A(n1199), .B(n1200), .C(n1203), .D(n1204), .S0(n1276), .S1(
        n1289), .Y(round_key[120]) );
  MXI4X1 U4686 ( .A(\key_mem[4][120] ), .B(\key_mem[5][120] ), .C(
        \key_mem[6][120] ), .D(\key_mem[7][120] ), .S0(n1390), .S1(n1332), .Y(
        n1203) );
  MXI3X1 U4687 ( .A(\key_mem[12][120] ), .B(\key_mem[13][120] ), .C(n1196), 
        .S0(n1380), .S1(n1334), .Y(n1204) );
  MXI4X1 U4688 ( .A(\key_mem[0][120] ), .B(\key_mem[1][120] ), .C(
        \key_mem[2][120] ), .D(\key_mem[3][120] ), .S0(n1390), .S1(n1333), .Y(
        n1199) );
  MXI4X1 U4689 ( .A(n1261), .B(n1262), .C(n1263), .D(n1264), .S0(n1276), .S1(
        n1289), .Y(round_key[127]) );
  MXI4X1 U4690 ( .A(\key_mem[4][127] ), .B(\key_mem[5][127] ), .C(
        \key_mem[6][127] ), .D(\key_mem[7][127] ), .S0(n1366), .S1(n1327), .Y(
        n1263) );
  MXI3X1 U4691 ( .A(\key_mem[12][127] ), .B(\key_mem[13][127] ), .C(n1260), 
        .S0(n1376), .S1(n1335), .Y(n1264) );
  MXI4X1 U4692 ( .A(\key_mem[0][127] ), .B(\key_mem[1][127] ), .C(
        \key_mem[2][127] ), .D(\key_mem[3][127] ), .S0(n1402), .S1(n1327), .Y(
        n1261) );
  MXI4X1 U4693 ( .A(n585), .B(n586), .C(n587), .D(n588), .S0(n1267), .S1(n1290), .Y(round_key[94]) );
  MXI4X1 U4694 ( .A(\key_mem[4][94] ), .B(\key_mem[5][94] ), .C(
        \key_mem[6][94] ), .D(\key_mem[7][94] ), .S0(n1398), .S1(n1326), .Y(
        n587) );
  MXI3X1 U4695 ( .A(\key_mem[12][94] ), .B(\key_mem[13][94] ), .C(n584), .S0(
        n1372), .S1(n1346), .Y(n588) );
  MXI4X1 U4696 ( .A(\key_mem[0][94] ), .B(\key_mem[1][94] ), .C(
        \key_mem[2][94] ), .D(\key_mem[3][94] ), .S0(n1398), .S1(n1326), .Y(
        n585) );
  MXI4X1 U4697 ( .A(n580), .B(n581), .C(n582), .D(n583), .S0(n1267), .S1(n1280), .Y(round_key[93]) );
  MXI4X1 U4698 ( .A(\key_mem[4][93] ), .B(\key_mem[5][93] ), .C(
        \key_mem[6][93] ), .D(\key_mem[7][93] ), .S0(n1398), .S1(n1326), .Y(
        n582) );
  MXI3X1 U4699 ( .A(\key_mem[12][93] ), .B(\key_mem[13][93] ), .C(n579), .S0(
        n1372), .S1(n1346), .Y(n583) );
  MXI4X1 U4700 ( .A(\key_mem[0][93] ), .B(\key_mem[1][93] ), .C(
        \key_mem[2][93] ), .D(\key_mem[3][93] ), .S0(n1398), .S1(n1326), .Y(
        n580) );
  MXI4X1 U4701 ( .A(n575), .B(n576), .C(n577), .D(n578), .S0(n1277), .S1(n1291), .Y(round_key[92]) );
  MXI4X1 U4702 ( .A(\key_mem[4][92] ), .B(\key_mem[5][92] ), .C(
        \key_mem[6][92] ), .D(\key_mem[7][92] ), .S0(n1399), .S1(n1326), .Y(
        n577) );
  MXI3X1 U4703 ( .A(\key_mem[12][92] ), .B(\key_mem[13][92] ), .C(n574), .S0(
        n1371), .S1(n1345), .Y(n578) );
  MXI4X1 U4704 ( .A(\key_mem[0][92] ), .B(\key_mem[1][92] ), .C(
        \key_mem[2][92] ), .D(\key_mem[3][92] ), .S0(n1399), .S1(n1326), .Y(
        n575) );
  MXI4X1 U4705 ( .A(n570), .B(n571), .C(n572), .D(n573), .S0(n1269), .S1(n1281), .Y(round_key[91]) );
  MXI4X1 U4706 ( .A(\key_mem[4][91] ), .B(\key_mem[5][91] ), .C(
        \key_mem[6][91] ), .D(\key_mem[7][91] ), .S0(n1399), .S1(n1325), .Y(
        n572) );
  MXI3X1 U4707 ( .A(\key_mem[12][91] ), .B(\key_mem[13][91] ), .C(n569), .S0(
        n1371), .S1(n1345), .Y(n573) );
  MXI4X1 U4708 ( .A(\key_mem[0][91] ), .B(\key_mem[1][91] ), .C(
        \key_mem[2][91] ), .D(\key_mem[3][91] ), .S0(n1399), .S1(n1325), .Y(
        n570) );
  MXI4X1 U4709 ( .A(n565), .B(n566), .C(n567), .D(n568), .S0(n1269), .S1(n1290), .Y(round_key[90]) );
  MXI4X1 U4710 ( .A(\key_mem[4][90] ), .B(\key_mem[5][90] ), .C(
        \key_mem[6][90] ), .D(\key_mem[7][90] ), .S0(n1399), .S1(n1325), .Y(
        n567) );
  MXI3X1 U4711 ( .A(\key_mem[12][90] ), .B(\key_mem[13][90] ), .C(n564), .S0(
        n1371), .S1(n1345), .Y(n568) );
  MXI4X1 U4712 ( .A(\key_mem[0][90] ), .B(\key_mem[1][90] ), .C(
        \key_mem[2][90] ), .D(\key_mem[3][90] ), .S0(n1399), .S1(n1325), .Y(
        n565) );
  MXI4X1 U4713 ( .A(n560), .B(n561), .C(n562), .D(n563), .S0(n1277), .S1(n1291), .Y(round_key[89]) );
  MXI3X1 U4714 ( .A(\key_mem[12][89] ), .B(\key_mem[13][89] ), .C(n559), .S0(
        n1370), .S1(n1345), .Y(n563) );
  MXI4X1 U4715 ( .A(\key_mem[4][89] ), .B(\key_mem[5][89] ), .C(
        \key_mem[6][89] ), .D(\key_mem[7][89] ), .S0(n1400), .S1(n1324), .Y(
        n562) );
  MXI4X1 U4716 ( .A(\key_mem[0][89] ), .B(\key_mem[1][89] ), .C(
        \key_mem[2][89] ), .D(\key_mem[3][89] ), .S0(n1399), .S1(n1325), .Y(
        n560) );
  MXI4X1 U4717 ( .A(n555), .B(n556), .C(n557), .D(n558), .S0(n1265), .S1(n1282), .Y(round_key[88]) );
  MXI3X1 U4718 ( .A(\key_mem[12][88] ), .B(\key_mem[13][88] ), .C(n554), .S0(
        n1370), .S1(n1345), .Y(n558) );
  MXI4X1 U4719 ( .A(\key_mem[4][88] ), .B(\key_mem[5][88] ), .C(
        \key_mem[6][88] ), .D(\key_mem[7][88] ), .S0(n1400), .S1(n1324), .Y(
        n557) );
  MXI4X1 U4720 ( .A(\key_mem[0][88] ), .B(\key_mem[1][88] ), .C(
        \key_mem[2][88] ), .D(\key_mem[3][88] ), .S0(n1400), .S1(n1324), .Y(
        n555) );
  MXI4X1 U4721 ( .A(n430), .B(n431), .C(n432), .D(n433), .S0(n1277), .S1(n1291), .Y(round_key[63]) );
  MXI4X1 U4722 ( .A(\key_mem[4][63] ), .B(\key_mem[5][63] ), .C(
        \key_mem[6][63] ), .D(\key_mem[7][63] ), .S0(n1386), .S1(n1315), .Y(
        n432) );
  MXI3X1 U4723 ( .A(\key_mem[12][63] ), .B(\key_mem[13][63] ), .C(n429), .S0(
        n1378), .S1(n1343), .Y(n433) );
  MXI4X1 U4724 ( .A(\key_mem[0][63] ), .B(\key_mem[1][63] ), .C(
        \key_mem[2][63] ), .D(\key_mem[3][63] ), .S0(n1386), .S1(n1315), .Y(
        n430) );
  MXI4X1 U4725 ( .A(n425), .B(n426), .C(n427), .D(n428), .S0(n1267), .S1(n1279), .Y(round_key[62]) );
  MXI4X1 U4726 ( .A(\key_mem[4][62] ), .B(\key_mem[5][62] ), .C(
        \key_mem[6][62] ), .D(\key_mem[7][62] ), .S0(n1385), .S1(n1314), .Y(
        n427) );
  MXI3X1 U4727 ( .A(\key_mem[12][62] ), .B(\key_mem[13][62] ), .C(n424), .S0(
        n1379), .S1(n1342), .Y(n428) );
  MXI4X1 U4728 ( .A(\key_mem[0][62] ), .B(\key_mem[1][62] ), .C(
        \key_mem[2][62] ), .D(\key_mem[3][62] ), .S0(n1386), .S1(n1314), .Y(
        n425) );
  MXI4X1 U4729 ( .A(n226), .B(n227), .C(n228), .D(n229), .S0(n1270), .S1(n1285), .Y(round_key[25]) );
  MXI3X1 U4730 ( .A(\key_mem[12][25] ), .B(\key_mem[13][25] ), .C(n225), .S0(
        n1370), .S1(n1339), .Y(n229) );
  MXI4X1 U4731 ( .A(\key_mem[4][25] ), .B(\key_mem[5][25] ), .C(
        \key_mem[6][25] ), .D(\key_mem[7][25] ), .S0(n1410), .S1(n1297), .Y(
        n228) );
  MXI4X1 U4732 ( .A(\key_mem[0][25] ), .B(\key_mem[1][25] ), .C(
        \key_mem[2][25] ), .D(\key_mem[3][25] ), .S0(n1410), .S1(n1305), .Y(
        n226) );
  MXI4X1 U4733 ( .A(n410), .B(n411), .C(n412), .D(n413), .S0(n1268), .S1(n1280), .Y(round_key[59]) );
  MXI4X1 U4734 ( .A(\key_mem[4][59] ), .B(\key_mem[5][59] ), .C(
        \key_mem[6][59] ), .D(\key_mem[7][59] ), .S0(n1383), .S1(n1313), .Y(
        n412) );
  MXI3X1 U4735 ( .A(\key_mem[12][59] ), .B(\key_mem[13][59] ), .C(n409), .S0(
        n1378), .S1(n1342), .Y(n413) );
  MXI4X1 U4736 ( .A(\key_mem[0][59] ), .B(\key_mem[1][59] ), .C(
        \key_mem[2][59] ), .D(\key_mem[3][59] ), .S0(n1384), .S1(n1313), .Y(
        n410) );
  MXI4X1 U4737 ( .A(n405), .B(n406), .C(n407), .D(n408), .S0(n1277), .S1(n1291), .Y(round_key[58]) );
  MXI4X1 U4738 ( .A(\key_mem[4][58] ), .B(\key_mem[5][58] ), .C(
        \key_mem[6][58] ), .D(\key_mem[7][58] ), .S0(n1383), .S1(n1313), .Y(
        n407) );
  MXI3X1 U4739 ( .A(\key_mem[12][58] ), .B(\key_mem[13][58] ), .C(n404), .S0(
        n1380), .S1(n1342), .Y(n408) );
  MXI4X1 U4740 ( .A(\key_mem[0][58] ), .B(\key_mem[1][58] ), .C(
        \key_mem[2][58] ), .D(\key_mem[3][58] ), .S0(n1383), .S1(n1313), .Y(
        n405) );
  MXI4X1 U4741 ( .A(n1239), .B(n1240), .C(n1243), .D(n1244), .S0(n1276), .S1(
        n1289), .Y(round_key[124]) );
  MXI4X1 U4742 ( .A(\key_mem[4][124] ), .B(\key_mem[5][124] ), .C(
        \key_mem[6][124] ), .D(\key_mem[7][124] ), .S0(n1389), .S1(n1329), .Y(
        n1243) );
  MXI3X1 U4743 ( .A(\key_mem[12][124] ), .B(\key_mem[13][124] ), .C(n1236), 
        .S0(n1377), .S1(n1334), .Y(n1244) );
  MXI4X1 U4744 ( .A(\key_mem[0][124] ), .B(\key_mem[1][124] ), .C(
        \key_mem[2][124] ), .D(\key_mem[3][124] ), .S0(n1389), .S1(n1329), .Y(
        n1239) );
  MXI4X1 U4745 ( .A(n1228), .B(n1231), .C(n1232), .D(n1235), .S0(n1276), .S1(
        n1289), .Y(round_key[123]) );
  MXI4X1 U4746 ( .A(\key_mem[4][123] ), .B(\key_mem[5][123] ), .C(
        \key_mem[6][123] ), .D(\key_mem[7][123] ), .S0(n1389), .S1(n1330), .Y(
        n1232) );
  MXI3X1 U4747 ( .A(\key_mem[12][123] ), .B(\key_mem[13][123] ), .C(n1227), 
        .S0(n1378), .S1(n1336), .Y(n1235) );
  MXI4X1 U4748 ( .A(\key_mem[0][123] ), .B(\key_mem[1][123] ), .C(
        \key_mem[2][123] ), .D(\key_mem[3][123] ), .S0(n1389), .S1(n1330), .Y(
        n1228) );
  MXI4X1 U4749 ( .A(n1219), .B(n1220), .C(n1223), .D(n1224), .S0(n1276), .S1(
        n1289), .Y(round_key[122]) );
  MXI4X1 U4750 ( .A(\key_mem[4][122] ), .B(\key_mem[5][122] ), .C(
        \key_mem[6][122] ), .D(\key_mem[7][122] ), .S0(n1390), .S1(n1295), .Y(
        n1223) );
  MXI3X1 U4751 ( .A(\key_mem[12][122] ), .B(\key_mem[13][122] ), .C(n1216), 
        .S0(n1378), .S1(n1336), .Y(n1224) );
  MXI4X1 U4752 ( .A(\key_mem[0][122] ), .B(\key_mem[1][122] ), .C(
        \key_mem[2][122] ), .D(\key_mem[3][122] ), .S0(n1389), .S1(n1295), .Y(
        n1219) );
  MXI4X1 U4753 ( .A(n592), .B(n721), .C(n744), .D(n745), .S0(n1266), .S1(n1291), .Y(round_key[95]) );
  MXI4X1 U4754 ( .A(\key_mem[4][95] ), .B(\key_mem[5][95] ), .C(
        \key_mem[6][95] ), .D(\key_mem[7][95] ), .S0(n1398), .S1(n1347), .Y(
        n744) );
  MXI3X1 U4755 ( .A(\key_mem[12][95] ), .B(\key_mem[13][95] ), .C(n589), .S0(
        n1373), .S1(n1346), .Y(n745) );
  MXI4X1 U4756 ( .A(\key_mem[0][95] ), .B(\key_mem[1][95] ), .C(
        \key_mem[2][95] ), .D(\key_mem[3][95] ), .S0(n1398), .S1(n1295), .Y(
        n592) );
  MXI4X1 U4757 ( .A(n1188), .B(n1191), .C(n1192), .D(n1195), .S0(n1276), .S1(
        n1289), .Y(round_key[119]) );
  MXI4X1 U4758 ( .A(\key_mem[4][119] ), .B(\key_mem[5][119] ), .C(
        \key_mem[6][119] ), .D(\key_mem[7][119] ), .S0(n1390), .S1(n1332), .Y(
        n1192) );
  MXI3X1 U4759 ( .A(\key_mem[12][119] ), .B(\key_mem[13][119] ), .C(n1187), 
        .S0(n1380), .S1(n1334), .Y(n1195) );
  MXI4X1 U4760 ( .A(\key_mem[0][119] ), .B(\key_mem[1][119] ), .C(
        \key_mem[2][119] ), .D(\key_mem[3][119] ), .S0(n1390), .S1(n1332), .Y(
        n1188) );
  MXI4X1 U4761 ( .A(n1155), .B(n1159), .C(n1163), .D(n1164), .S0(n1275), .S1(
        n1280), .Y(round_key[116]) );
  MXI4X1 U4762 ( .A(\key_mem[4][116] ), .B(\key_mem[5][116] ), .C(
        \key_mem[6][116] ), .D(\key_mem[7][116] ), .S0(n1391), .S1(n1297), .Y(
        n1163) );
  MXI3X1 U4763 ( .A(\key_mem[12][116] ), .B(\key_mem[13][116] ), .C(n1151), 
        .S0(n1380), .S1(n1336), .Y(n1164) );
  MXI4X1 U4764 ( .A(\key_mem[0][116] ), .B(\key_mem[1][116] ), .C(
        \key_mem[2][116] ), .D(\key_mem[3][116] ), .S0(n1391), .S1(n1301), .Y(
        n1155) );
  MXI4X1 U4765 ( .A(n535), .B(n536), .C(n537), .D(n538), .S0(n1278), .S1(n1292), .Y(round_key[84]) );
  MXI3X1 U4766 ( .A(\key_mem[12][84] ), .B(\key_mem[13][84] ), .C(n534), .S0(
        n1352), .S1(n1345), .Y(n538) );
  MXI4X1 U4767 ( .A(\key_mem[4][84] ), .B(\key_mem[5][84] ), .C(
        \key_mem[6][84] ), .D(\key_mem[7][84] ), .S0(n1401), .S1(n1323), .Y(
        n537) );
  MXI4X1 U4768 ( .A(\key_mem[0][84] ), .B(\key_mem[1][84] ), .C(
        \key_mem[2][84] ), .D(\key_mem[3][84] ), .S0(n1401), .S1(n1323), .Y(
        n535) );
  MXI4X1 U4769 ( .A(n1135), .B(n1139), .C(n1143), .D(n1147), .S0(n1275), .S1(
        N33), .Y(round_key[115]) );
  MXI4X1 U4770 ( .A(\key_mem[4][115] ), .B(\key_mem[5][115] ), .C(
        \key_mem[6][115] ), .D(\key_mem[7][115] ), .S0(n1392), .S1(n1308), .Y(
        n1143) );
  MXI3X1 U4771 ( .A(\key_mem[12][115] ), .B(\key_mem[13][115] ), .C(n1132), 
        .S0(n1378), .S1(n1336), .Y(n1147) );
  MXI4X1 U4772 ( .A(\key_mem[0][115] ), .B(\key_mem[1][115] ), .C(
        \key_mem[2][115] ), .D(\key_mem[3][115] ), .S0(n1392), .S1(n1294), .Y(
        n1135) );
  MXI4X1 U4773 ( .A(n1124), .B(n1125), .C(n1128), .D(n1131), .S0(n1275), .S1(
        n1292), .Y(round_key[114]) );
  MXI4X1 U4774 ( .A(\key_mem[4][114] ), .B(\key_mem[5][114] ), .C(
        \key_mem[6][114] ), .D(\key_mem[7][114] ), .S0(n1392), .S1(n1311), .Y(
        n1128) );
  MXI3X1 U4775 ( .A(\key_mem[12][114] ), .B(\key_mem[13][114] ), .C(n1120), 
        .S0(n1379), .S1(n1335), .Y(n1131) );
  MXI4X1 U4776 ( .A(\key_mem[0][114] ), .B(\key_mem[1][114] ), .C(
        \key_mem[2][114] ), .D(\key_mem[3][114] ), .S0(n1392), .S1(n1310), .Y(
        n1124) );
  MXI4X1 U4777 ( .A(n525), .B(n526), .C(n527), .D(n528), .S0(n1269), .S1(n1279), .Y(round_key[82]) );
  MXI3X1 U4778 ( .A(\key_mem[12][82] ), .B(\key_mem[13][82] ), .C(n524), .S0(
        n1369), .S1(n1344), .Y(n528) );
  MXI4X1 U4779 ( .A(\key_mem[4][82] ), .B(\key_mem[5][82] ), .C(
        \key_mem[6][82] ), .D(\key_mem[7][82] ), .S0(n1402), .S1(n1322), .Y(
        n527) );
  MXI4X1 U4780 ( .A(\key_mem[0][82] ), .B(\key_mem[1][82] ), .C(
        \key_mem[2][82] ), .D(\key_mem[3][82] ), .S0(n1402), .S1(n1322), .Y(
        n525) );
  MXI4X1 U4781 ( .A(n167), .B(n168), .C(n169), .D(n170), .S0(n1270), .S1(n1285), .Y(round_key[18]) );
  MXI3X1 U4782 ( .A(\key_mem[12][18] ), .B(\key_mem[13][18] ), .C(n166), .S0(
        n1369), .S1(n1338), .Y(n170) );
  MXI4X1 U4783 ( .A(\key_mem[4][18] ), .B(\key_mem[5][18] ), .C(
        \key_mem[6][18] ), .D(\key_mem[7][18] ), .S0(n1408), .S1(n1302), .Y(
        n169) );
  MXI4X1 U4784 ( .A(\key_mem[0][18] ), .B(\key_mem[1][18] ), .C(
        \key_mem[2][18] ), .D(\key_mem[3][18] ), .S0(n1408), .S1(n1303), .Y(
        n167) );
  MXI4X1 U4785 ( .A(n520), .B(n521), .C(n522), .D(n523), .S0(n1268), .S1(N33), 
        .Y(round_key[81]) );
  MXI4X1 U4786 ( .A(\key_mem[4][81] ), .B(\key_mem[5][81] ), .C(
        \key_mem[6][81] ), .D(\key_mem[7][81] ), .S0(n1402), .S1(n1321), .Y(
        n522) );
  MXI3X1 U4787 ( .A(\key_mem[12][81] ), .B(\key_mem[13][81] ), .C(n519), .S0(
        n1376), .S1(n1344), .Y(n523) );
  MXI4X1 U4788 ( .A(\key_mem[0][81] ), .B(\key_mem[1][81] ), .C(
        \key_mem[2][81] ), .D(\key_mem[3][81] ), .S0(n1402), .S1(n1322), .Y(
        n520) );
  MXI4X1 U4789 ( .A(n162), .B(n163), .C(n164), .D(n165), .S0(n1278), .S1(n1284), .Y(round_key[17]) );
  MXI3X1 U4790 ( .A(\key_mem[12][17] ), .B(\key_mem[13][17] ), .C(n161), .S0(
        n1369), .S1(n1338), .Y(n165) );
  MXI4X1 U4791 ( .A(\key_mem[4][17] ), .B(\key_mem[5][17] ), .C(
        \key_mem[6][17] ), .D(\key_mem[7][17] ), .S0(n1407), .S1(n1293), .Y(
        n164) );
  MXI4X1 U4792 ( .A(\key_mem[0][17] ), .B(\key_mem[1][17] ), .C(
        \key_mem[2][17] ), .D(\key_mem[3][17] ), .S0(n1408), .S1(n1308), .Y(
        n162) );
  MXI4X1 U4793 ( .A(n1104), .B(n1108), .C(n1112), .D(n1116), .S0(n1275), .S1(
        N33), .Y(round_key[113]) );
  MXI4X1 U4794 ( .A(\key_mem[4][113] ), .B(\key_mem[5][113] ), .C(
        \key_mem[6][113] ), .D(\key_mem[7][113] ), .S0(n1392), .S1(n1312), .Y(
        n1112) );
  MXI3X1 U4795 ( .A(\key_mem[12][113] ), .B(\key_mem[13][113] ), .C(n1100), 
        .S0(n1378), .S1(n1335), .Y(n1116) );
  MXI4X1 U4796 ( .A(\key_mem[0][113] ), .B(\key_mem[1][113] ), .C(
        \key_mem[2][113] ), .D(\key_mem[3][113] ), .S0(n1392), .S1(n1312), .Y(
        n1104) );
  MXI4X1 U4797 ( .A(n515), .B(n516), .C(n517), .D(n518), .S0(n1268), .S1(n1279), .Y(round_key[80]) );
  MXI3X1 U4798 ( .A(\key_mem[12][80] ), .B(\key_mem[13][80] ), .C(n514), .S0(
        n1369), .S1(n1344), .Y(n518) );
  MXI4X1 U4799 ( .A(\key_mem[4][80] ), .B(\key_mem[5][80] ), .C(
        \key_mem[6][80] ), .D(\key_mem[7][80] ), .S0(n1381), .S1(n1321), .Y(
        n517) );
  MXI4X1 U4800 ( .A(\key_mem[0][80] ), .B(\key_mem[1][80] ), .C(
        \key_mem[2][80] ), .D(\key_mem[3][80] ), .S0(n1395), .S1(n1321), .Y(
        n515) );
  MXI4X1 U4801 ( .A(n216), .B(n217), .C(n218), .D(n219), .S0(n1270), .S1(n1285), .Y(round_key[23]) );
  MXI3X1 U4802 ( .A(\key_mem[12][23] ), .B(\key_mem[13][23] ), .C(n215), .S0(
        n1353), .S1(n1338), .Y(n219) );
  MXI4X1 U4803 ( .A(\key_mem[4][23] ), .B(\key_mem[5][23] ), .C(
        \key_mem[6][23] ), .D(\key_mem[7][23] ), .S0(n1409), .S1(n1304), .Y(
        n218) );
  MXI4X1 U4804 ( .A(\key_mem[0][23] ), .B(\key_mem[1][23] ), .C(
        \key_mem[2][23] ), .D(\key_mem[3][23] ), .S0(n1409), .S1(n1298), .Y(
        n216) );
  MXI4X1 U4805 ( .A(n1179), .B(n1180), .C(n1183), .D(n1184), .S0(n1276), .S1(
        n1289), .Y(round_key[118]) );
  MXI4X1 U4806 ( .A(\key_mem[4][118] ), .B(\key_mem[5][118] ), .C(
        \key_mem[6][118] ), .D(\key_mem[7][118] ), .S0(n1391), .S1(n1309), .Y(
        n1183) );
  MXI3X1 U4807 ( .A(\key_mem[12][118] ), .B(\key_mem[13][118] ), .C(n1176), 
        .S0(n1379), .S1(n1335), .Y(n1184) );
  MXI4X1 U4808 ( .A(\key_mem[0][118] ), .B(\key_mem[1][118] ), .C(
        \key_mem[2][118] ), .D(\key_mem[3][118] ), .S0(n1391), .S1(n1309), .Y(
        n1179) );
  MXI4X1 U4809 ( .A(n540), .B(n541), .C(n542), .D(n543), .S0(n1266), .S1(n1279), .Y(round_key[85]) );
  MXI3X1 U4810 ( .A(\key_mem[12][85] ), .B(\key_mem[13][85] ), .C(n539), .S0(
        n1352), .S1(n1345), .Y(n543) );
  MXI4X1 U4811 ( .A(\key_mem[4][85] ), .B(\key_mem[5][85] ), .C(
        \key_mem[6][85] ), .D(\key_mem[7][85] ), .S0(n1401), .S1(n1323), .Y(
        n542) );
  MXI4X1 U4812 ( .A(\key_mem[0][85] ), .B(\key_mem[1][85] ), .C(
        \key_mem[2][85] ), .D(\key_mem[3][85] ), .S0(n1401), .S1(n1323), .Y(
        n540) );
  MXI4X1 U4813 ( .A(n380), .B(n381), .C(n382), .D(n383), .S0(n1273), .S1(n1288), .Y(round_key[53]) );
  MXI4X1 U4814 ( .A(\key_mem[4][53] ), .B(\key_mem[5][53] ), .C(
        \key_mem[6][53] ), .D(\key_mem[7][53] ), .S0(n1411), .S1(n1311), .Y(
        n382) );
  MXI3X1 U4815 ( .A(\key_mem[12][53] ), .B(\key_mem[13][53] ), .C(n379), .S0(
        n1376), .S1(n1342), .Y(n383) );
  MXI4X1 U4816 ( .A(\key_mem[0][53] ), .B(\key_mem[1][53] ), .C(
        \key_mem[2][53] ), .D(\key_mem[3][53] ), .S0(n1411), .S1(n1311), .Y(
        n380) );
  MXI4X1 U4817 ( .A(n157), .B(n158), .C(n159), .D(n160), .S0(n1265), .S1(n1284), .Y(round_key[16]) );
  MXI3X1 U4818 ( .A(\key_mem[12][16] ), .B(\key_mem[13][16] ), .C(n156), .S0(
        n1369), .S1(n1338), .Y(n160) );
  MXI4X1 U4819 ( .A(\key_mem[4][16] ), .B(\key_mem[5][16] ), .C(
        \key_mem[6][16] ), .D(\key_mem[7][16] ), .S0(n1407), .S1(n1330), .Y(
        n159) );
  MXI4X1 U4820 ( .A(\key_mem[0][16] ), .B(\key_mem[1][16] ), .C(
        \key_mem[2][16] ), .D(\key_mem[3][16] ), .S0(n1407), .S1(n1330), .Y(
        n157) );
  MXI4X1 U4821 ( .A(n1168), .B(n1171), .C(n1172), .D(n1175), .S0(n1275), .S1(
        n1279), .Y(round_key[117]) );
  MXI4X1 U4822 ( .A(\key_mem[4][117] ), .B(\key_mem[5][117] ), .C(
        \key_mem[6][117] ), .D(\key_mem[7][117] ), .S0(n1391), .S1(n1348), .Y(
        n1172) );
  MXI3X1 U4823 ( .A(\key_mem[12][117] ), .B(\key_mem[13][117] ), .C(n1167), 
        .S0(n1379), .S1(n1334), .Y(n1175) );
  MXI4X1 U4824 ( .A(\key_mem[0][117] ), .B(\key_mem[1][117] ), .C(
        \key_mem[2][117] ), .D(\key_mem[3][117] ), .S0(n1391), .S1(n1348), .Y(
        n1168) );
  MXI4X1 U4825 ( .A(n340), .B(n341), .C(n342), .D(n343), .S0(n1272), .S1(n1287), .Y(round_key[45]) );
  MXI4X1 U4826 ( .A(\key_mem[4][45] ), .B(\key_mem[5][45] ), .C(
        \key_mem[6][45] ), .D(\key_mem[7][45] ), .S0(n1413), .S1(n1302), .Y(
        n342) );
  MXI3X1 U4827 ( .A(\key_mem[12][45] ), .B(\key_mem[13][45] ), .C(n339), .S0(
        n1376), .S1(n1341), .Y(n343) );
  MXI4X1 U4828 ( .A(\key_mem[0][45] ), .B(\key_mem[1][45] ), .C(
        \key_mem[2][45] ), .D(\key_mem[3][45] ), .S0(n1413), .S1(n1297), .Y(
        n340) );
  MXI4X1 U4829 ( .A(n1023), .B(n1027), .C(n1031), .D(n1036), .S0(n1275), .S1(
        n1291), .Y(round_key[109]) );
  MXI4X1 U4830 ( .A(\key_mem[4][109] ), .B(\key_mem[5][109] ), .C(
        \key_mem[6][109] ), .D(\key_mem[7][109] ), .S0(n1393), .S1(n1318), .Y(
        n1031) );
  MXI3X1 U4831 ( .A(\key_mem[12][109] ), .B(\key_mem[13][109] ), .C(n1019), 
        .S0(n1376), .S1(n1336), .Y(n1036) );
  MXI4X1 U4832 ( .A(\key_mem[0][109] ), .B(\key_mem[1][109] ), .C(
        \key_mem[2][109] ), .D(\key_mem[3][109] ), .S0(n1393), .S1(n1318), .Y(
        n1023) );
  MXI4X1 U4833 ( .A(n385), .B(n386), .C(n387), .D(n388), .S0(n1273), .S1(n1288), .Y(round_key[54]) );
  MXI4X1 U4834 ( .A(\key_mem[4][54] ), .B(\key_mem[5][54] ), .C(
        \key_mem[6][54] ), .D(\key_mem[7][54] ), .S0(n1410), .S1(n1311), .Y(
        n387) );
  MXI3X1 U4835 ( .A(\key_mem[12][54] ), .B(\key_mem[13][54] ), .C(n384), .S0(
        n1376), .S1(n1342), .Y(n388) );
  MXI4X1 U4836 ( .A(\key_mem[0][54] ), .B(\key_mem[1][54] ), .C(
        \key_mem[2][54] ), .D(\key_mem[3][54] ), .S0(n1385), .S1(n1311), .Y(
        n385) );
  MXI4X1 U4837 ( .A(n1044), .B(n1048), .C(n1052), .D(n1056), .S0(n1275), .S1(
        n1282), .Y(round_key[110]) );
  MXI4X1 U4838 ( .A(\key_mem[4][110] ), .B(\key_mem[5][110] ), .C(
        \key_mem[6][110] ), .D(\key_mem[7][110] ), .S0(n1393), .S1(n1317), .Y(
        n1052) );
  MXI3X1 U4839 ( .A(\key_mem[12][110] ), .B(\key_mem[13][110] ), .C(n1040), 
        .S0(n1377), .S1(n1335), .Y(n1056) );
  MXI4X1 U4840 ( .A(\key_mem[0][110] ), .B(\key_mem[1][110] ), .C(
        \key_mem[2][110] ), .D(\key_mem[3][110] ), .S0(n1393), .S1(n1316), .Y(
        n1044) );
  MXI4X1 U4841 ( .A(n345), .B(n346), .C(n347), .D(n348), .S0(n1272), .S1(n1287), .Y(round_key[46]) );
  MXI4X1 U4842 ( .A(\key_mem[4][46] ), .B(\key_mem[5][46] ), .C(
        \key_mem[6][46] ), .D(\key_mem[7][46] ), .S0(n1413), .S1(n1306), .Y(
        n347) );
  MXI3X1 U4843 ( .A(\key_mem[12][46] ), .B(\key_mem[13][46] ), .C(n344), .S0(
        n1377), .S1(n1341), .Y(n348) );
  MXI4X1 U4844 ( .A(\key_mem[0][46] ), .B(\key_mem[1][46] ), .C(
        \key_mem[2][46] ), .D(\key_mem[3][46] ), .S0(n1413), .S1(n1299), .Y(
        n345) );
  MXI4X1 U4845 ( .A(n211), .B(n212), .C(n213), .D(n214), .S0(n1270), .S1(n1285), .Y(round_key[22]) );
  MXI3X1 U4846 ( .A(\key_mem[12][22] ), .B(\key_mem[13][22] ), .C(n210), .S0(
        N31), .S1(n1338), .Y(n214) );
  MXI4X1 U4847 ( .A(\key_mem[4][22] ), .B(\key_mem[5][22] ), .C(
        \key_mem[6][22] ), .D(\key_mem[7][22] ), .S0(n1409), .S1(n1305), .Y(
        n213) );
  MXI4X1 U4848 ( .A(\key_mem[0][22] ), .B(\key_mem[1][22] ), .C(
        \key_mem[2][22] ), .D(\key_mem[3][22] ), .S0(n1409), .S1(n1296), .Y(
        n211) );
  MXI4X1 U4849 ( .A(n505), .B(n506), .C(n507), .D(n508), .S0(n1277), .S1(n1281), .Y(round_key[78]) );
  MXI3X1 U4850 ( .A(\key_mem[12][78] ), .B(\key_mem[13][78] ), .C(n504), .S0(
        n1352), .S1(n1344), .Y(n508) );
  MXI4X1 U4851 ( .A(\key_mem[4][78] ), .B(\key_mem[5][78] ), .C(
        \key_mem[6][78] ), .D(\key_mem[7][78] ), .S0(n1381), .S1(n1320), .Y(
        n507) );
  MXI4X1 U4852 ( .A(\key_mem[0][78] ), .B(\key_mem[1][78] ), .C(
        \key_mem[2][78] ), .D(\key_mem[3][78] ), .S0(n1382), .S1(n1320), .Y(
        n505) );
  MXI4X1 U4853 ( .A(n147), .B(n148), .C(n149), .D(n150), .S0(n1265), .S1(n1284), .Y(round_key[14]) );
  MXI3X1 U4854 ( .A(\key_mem[12][14] ), .B(\key_mem[13][14] ), .C(n146), .S0(
        n1356), .S1(n1338), .Y(n150) );
  MXI4X1 U4855 ( .A(\key_mem[4][14] ), .B(\key_mem[5][14] ), .C(
        \key_mem[6][14] ), .D(\key_mem[7][14] ), .S0(n1407), .S1(n1330), .Y(
        n149) );
  MXI4X1 U4856 ( .A(\key_mem[0][14] ), .B(\key_mem[1][14] ), .C(
        \key_mem[2][14] ), .D(\key_mem[3][14] ), .S0(n1407), .S1(n1330), .Y(
        n147) );
  MXI4X1 U4857 ( .A(n500), .B(n501), .C(n502), .D(n503), .S0(n1269), .S1(n1292), .Y(round_key[77]) );
  MXI3X1 U4858 ( .A(\key_mem[12][77] ), .B(\key_mem[13][77] ), .C(n499), .S0(
        n1370), .S1(n1344), .Y(n503) );
  MXI4X1 U4859 ( .A(\key_mem[4][77] ), .B(\key_mem[5][77] ), .C(
        \key_mem[6][77] ), .D(\key_mem[7][77] ), .S0(n1383), .S1(n1320), .Y(
        n502) );
  MXI4X1 U4860 ( .A(\key_mem[0][77] ), .B(\key_mem[1][77] ), .C(
        \key_mem[2][77] ), .D(\key_mem[3][77] ), .S0(n1382), .S1(n1320), .Y(
        n500) );
  MXI4X1 U4861 ( .A(n142), .B(n143), .C(n144), .D(n145), .S0(n1265), .S1(n1284), .Y(round_key[13]) );
  MXI3X1 U4862 ( .A(\key_mem[12][13] ), .B(\key_mem[13][13] ), .C(n141), .S0(
        n1350), .S1(n1337), .Y(n145) );
  MXI4X1 U4863 ( .A(\key_mem[4][13] ), .B(\key_mem[5][13] ), .C(
        \key_mem[6][13] ), .D(\key_mem[7][13] ), .S0(n1406), .S1(n1329), .Y(
        n144) );
  MXI4X1 U4864 ( .A(\key_mem[0][13] ), .B(\key_mem[1][13] ), .C(
        \key_mem[2][13] ), .D(\key_mem[3][13] ), .S0(n1406), .S1(n1329), .Y(
        n142) );
  MXI4X1 U4865 ( .A(n137), .B(n138), .C(n139), .D(n140), .S0(n1265), .S1(n1284), .Y(round_key[12]) );
  MXI3X1 U4866 ( .A(\key_mem[12][12] ), .B(\key_mem[13][12] ), .C(n136), .S0(
        n1351), .S1(n1337), .Y(n140) );
  MXI4X1 U4867 ( .A(\key_mem[4][12] ), .B(\key_mem[5][12] ), .C(
        \key_mem[6][12] ), .D(\key_mem[7][12] ), .S0(n1406), .S1(n1329), .Y(
        n139) );
  MXI4X1 U4868 ( .A(\key_mem[0][12] ), .B(\key_mem[1][12] ), .C(
        \key_mem[2][12] ), .D(\key_mem[3][12] ), .S0(n1406), .S1(n1329), .Y(
        n137) );
  MXI4X1 U4869 ( .A(n475), .B(n476), .C(n477), .D(n478), .S0(n1277), .S1(n1281), .Y(round_key[72]) );
  MXI4X1 U4870 ( .A(\key_mem[4][72] ), .B(\key_mem[5][72] ), .C(
        \key_mem[6][72] ), .D(\key_mem[7][72] ), .S0(n1385), .S1(n1318), .Y(
        n477) );
  MXI3X1 U4871 ( .A(\key_mem[12][72] ), .B(\key_mem[13][72] ), .C(n474), .S0(
        n1373), .S1(n1343), .Y(n478) );
  MXI4X1 U4872 ( .A(\key_mem[0][72] ), .B(\key_mem[1][72] ), .C(
        \key_mem[2][72] ), .D(\key_mem[3][72] ), .S0(n1385), .S1(n1318), .Y(
        n475) );
  MXI4X1 U4873 ( .A(n117), .B(n118), .C(n119), .D(n120), .S0(n1265), .S1(n1284), .Y(round_key[8]) );
  MXI4X1 U4874 ( .A(\key_mem[4][8] ), .B(\key_mem[5][8] ), .C(\key_mem[6][8] ), 
        .D(\key_mem[7][8] ), .S0(n1405), .S1(n1299), .Y(n119) );
  MXI3X1 U4875 ( .A(\key_mem[12][8] ), .B(\key_mem[13][8] ), .C(n116), .S0(
        n1371), .S1(n1337), .Y(n120) );
  MXI4X1 U4876 ( .A(\key_mem[0][8] ), .B(\key_mem[1][8] ), .C(\key_mem[2][8] ), 
        .D(\key_mem[3][8] ), .S0(n1405), .S1(n1303), .Y(n117) );
  MXI4X1 U4877 ( .A(n1084), .B(n1088), .C(n1092), .D(n1096), .S0(n1275), .S1(
        n1279), .Y(round_key[112]) );
  MXI4X1 U4878 ( .A(\key_mem[4][112] ), .B(\key_mem[5][112] ), .C(
        \key_mem[6][112] ), .D(\key_mem[7][112] ), .S0(n1393), .S1(n1314), .Y(
        n1092) );
  MXI3X1 U4879 ( .A(\key_mem[12][112] ), .B(\key_mem[13][112] ), .C(n1080), 
        .S0(n1378), .S1(n1334), .Y(n1096) );
  MXI4X1 U4880 ( .A(\key_mem[0][112] ), .B(\key_mem[1][112] ), .C(
        \key_mem[2][112] ), .D(\key_mem[3][112] ), .S0(n1392), .S1(n1313), .Y(
        n1084) );
  MXI4X1 U4881 ( .A(n350), .B(n351), .C(n352), .D(n353), .S0(n1272), .S1(n1287), .Y(round_key[47]) );
  MXI4X1 U4882 ( .A(\key_mem[4][47] ), .B(\key_mem[5][47] ), .C(
        \key_mem[6][47] ), .D(\key_mem[7][47] ), .S0(n1413), .S1(n1308), .Y(
        n352) );
  MXI3X1 U4883 ( .A(\key_mem[12][47] ), .B(\key_mem[13][47] ), .C(n349), .S0(
        n1380), .S1(n1341), .Y(n353) );
  MXI4X1 U4884 ( .A(\key_mem[0][47] ), .B(\key_mem[1][47] ), .C(
        \key_mem[2][47] ), .D(\key_mem[3][47] ), .S0(n1412), .S1(n1303), .Y(
        n350) );
  MXI4X1 U4885 ( .A(n470), .B(n471), .C(n472), .D(n473), .S0(n1277), .S1(n1279), .Y(round_key[71]) );
  MXI4X1 U4886 ( .A(\key_mem[4][71] ), .B(\key_mem[5][71] ), .C(
        \key_mem[6][71] ), .D(\key_mem[7][71] ), .S0(n1386), .S1(n1318), .Y(
        n472) );
  MXI3X1 U4887 ( .A(\key_mem[12][71] ), .B(\key_mem[13][71] ), .C(n469), .S0(
        n1373), .S1(n1343), .Y(n473) );
  MXI4X1 U4888 ( .A(\key_mem[0][71] ), .B(\key_mem[1][71] ), .C(
        \key_mem[2][71] ), .D(\key_mem[3][71] ), .S0(n1385), .S1(n1318), .Y(
        n470) );
  MXI4X1 U4889 ( .A(n152), .B(n153), .C(n154), .D(n155), .S0(n1269), .S1(n1284), .Y(round_key[15]) );
  MXI3X1 U4890 ( .A(\key_mem[12][15] ), .B(\key_mem[13][15] ), .C(n151), .S0(
        n1350), .S1(n1338), .Y(n155) );
  MXI4X1 U4891 ( .A(\key_mem[4][15] ), .B(\key_mem[5][15] ), .C(
        \key_mem[6][15] ), .D(\key_mem[7][15] ), .S0(n1407), .S1(n1330), .Y(
        n154) );
  MXI4X1 U4892 ( .A(\key_mem[0][15] ), .B(\key_mem[1][15] ), .C(
        \key_mem[2][15] ), .D(\key_mem[3][15] ), .S0(n1407), .S1(n1330), .Y(
        n152) );
  MXI4X1 U4893 ( .A(n310), .B(n311), .C(n312), .D(n313), .S0(n1272), .S1(n1287), .Y(round_key[39]) );
  MXI4X1 U4894 ( .A(\key_mem[4][39] ), .B(\key_mem[5][39] ), .C(
        \key_mem[6][39] ), .D(\key_mem[7][39] ), .S0(n1415), .S1(n1348), .Y(
        n312) );
  MXI3X1 U4895 ( .A(\key_mem[12][39] ), .B(\key_mem[13][39] ), .C(n309), .S0(
        n1375), .S1(n1340), .Y(n313) );
  MXI4X1 U4896 ( .A(\key_mem[0][39] ), .B(\key_mem[1][39] ), .C(
        \key_mem[2][39] ), .D(\key_mem[3][39] ), .S0(n1415), .S1(n1299), .Y(
        n310) );
  MXI4X1 U4897 ( .A(n1064), .B(n1068), .C(n1072), .D(n1076), .S0(n1275), .S1(
        n1291), .Y(round_key[111]) );
  MXI4X1 U4898 ( .A(\key_mem[4][111] ), .B(\key_mem[5][111] ), .C(
        \key_mem[6][111] ), .D(\key_mem[7][111] ), .S0(n1393), .S1(n1315), .Y(
        n1072) );
  MXI3X1 U4899 ( .A(\key_mem[12][111] ), .B(\key_mem[13][111] ), .C(n1060), 
        .S0(n1378), .S1(n1335), .Y(n1076) );
  MXI4X1 U4900 ( .A(\key_mem[0][111] ), .B(\key_mem[1][111] ), .C(
        \key_mem[2][111] ), .D(\key_mem[3][111] ), .S0(n1393), .S1(n1315), .Y(
        n1064) );
  MXI4X1 U4901 ( .A(n112), .B(n113), .C(n114), .D(n115), .S0(n1269), .S1(n1283), .Y(round_key[7]) );
  MXI4X1 U4902 ( .A(\key_mem[4][7] ), .B(\key_mem[5][7] ), .C(\key_mem[6][7] ), 
        .D(\key_mem[7][7] ), .S0(n1404), .S1(n1300), .Y(n114) );
  MXI3X1 U4903 ( .A(\key_mem[12][7] ), .B(\key_mem[13][7] ), .C(n111), .S0(
        n1371), .S1(n1337), .Y(n115) );
  MXI4X1 U4904 ( .A(\key_mem[0][7] ), .B(\key_mem[1][7] ), .C(\key_mem[2][7] ), 
        .D(\key_mem[3][7] ), .S0(n1405), .S1(n1306), .Y(n112) );
  MXI4X1 U4905 ( .A(n510), .B(n511), .C(n512), .D(n513), .S0(n1277), .S1(n1279), .Y(round_key[79]) );
  MXI4X1 U4906 ( .A(\key_mem[4][79] ), .B(\key_mem[5][79] ), .C(
        \key_mem[6][79] ), .D(\key_mem[7][79] ), .S0(n1380), .S1(n1321), .Y(
        n512) );
  MXI3X1 U4907 ( .A(\key_mem[12][79] ), .B(\key_mem[13][79] ), .C(n509), .S0(
        n1369), .S1(n1344), .Y(n513) );
  MXI4X1 U4908 ( .A(\key_mem[0][79] ), .B(\key_mem[1][79] ), .C(
        \key_mem[2][79] ), .D(\key_mem[3][79] ), .S0(n1381), .S1(n1321), .Y(
        n510) );
  MXI4X1 U4909 ( .A(n955), .B(n956), .C(n959), .D(n960), .S0(n1274), .S1(n1290), .Y(round_key[103]) );
  MXI4X1 U4910 ( .A(\key_mem[4][103] ), .B(\key_mem[5][103] ), .C(
        \key_mem[6][103] ), .D(\key_mem[7][103] ), .S0(n1395), .S1(n1348), .Y(
        n959) );
  MXI3X1 U4911 ( .A(\key_mem[12][103] ), .B(\key_mem[13][103] ), .C(n952), 
        .S0(n1375), .S1(n1336), .Y(n960) );
  MXI4X1 U4912 ( .A(\key_mem[0][103] ), .B(\key_mem[1][103] ), .C(
        \key_mem[2][103] ), .D(\key_mem[3][103] ), .S0(n1395), .S1(n1303), .Y(
        n955) );
  MXI4X1 U4913 ( .A(n305), .B(n306), .C(n307), .D(n308), .S0(n1272), .S1(n1287), .Y(round_key[38]) );
  MXI4X1 U4914 ( .A(\key_mem[4][38] ), .B(\key_mem[5][38] ), .C(
        \key_mem[6][38] ), .D(\key_mem[7][38] ), .S0(n1415), .S1(n1294), .Y(
        n307) );
  MXI3X1 U4915 ( .A(\key_mem[12][38] ), .B(\key_mem[13][38] ), .C(n304), .S0(
        n1375), .S1(n1340), .Y(n308) );
  MXI4X1 U4916 ( .A(\key_mem[0][38] ), .B(\key_mem[1][38] ), .C(
        \key_mem[2][38] ), .D(\key_mem[3][38] ), .S0(n1415), .S1(n1347), .Y(
        n305) );
  MXI4X1 U4917 ( .A(n465), .B(n466), .C(n467), .D(n468), .S0(n1266), .S1(n1281), .Y(round_key[70]) );
  MXI4X1 U4918 ( .A(\key_mem[4][70] ), .B(\key_mem[5][70] ), .C(
        \key_mem[6][70] ), .D(\key_mem[7][70] ), .S0(n1386), .S1(n1317), .Y(
        n467) );
  MXI3X1 U4919 ( .A(\key_mem[12][70] ), .B(\key_mem[13][70] ), .C(n464), .S0(
        n1374), .S1(n1343), .Y(n468) );
  MXI4X1 U4920 ( .A(\key_mem[0][70] ), .B(\key_mem[1][70] ), .C(
        \key_mem[2][70] ), .D(\key_mem[3][70] ), .S0(n1386), .S1(n1317), .Y(
        n465) );
  MXI4X1 U4921 ( .A(n944), .B(n947), .C(n948), .D(n951), .S0(n1274), .S1(n1290), .Y(round_key[102]) );
  MXI4X1 U4922 ( .A(\key_mem[4][102] ), .B(\key_mem[5][102] ), .C(
        \key_mem[6][102] ), .D(\key_mem[7][102] ), .S0(n1396), .S1(n1327), .Y(
        n948) );
  MXI3X1 U4923 ( .A(\key_mem[12][102] ), .B(\key_mem[13][102] ), .C(n943), 
        .S0(n1374), .S1(n1341), .Y(n951) );
  MXI4X1 U4924 ( .A(\key_mem[0][102] ), .B(\key_mem[1][102] ), .C(
        \key_mem[2][102] ), .D(\key_mem[3][102] ), .S0(n1396), .S1(n1347), .Y(
        n944) );
  MXI4X1 U4925 ( .A(n102), .B(n103), .C(n104), .D(n105), .S0(n1269), .S1(n1283), .Y(round_key[5]) );
  MXI4X1 U4926 ( .A(\key_mem[4][5] ), .B(\key_mem[5][5] ), .C(\key_mem[6][5] ), 
        .D(\key_mem[7][5] ), .S0(n1404), .S1(n1294), .Y(n104) );
  MXI3X1 U4927 ( .A(\key_mem[12][5] ), .B(\key_mem[13][5] ), .C(n101), .S0(
        n1371), .S1(n1337), .Y(n105) );
  MXI4X1 U4928 ( .A(\key_mem[0][5] ), .B(\key_mem[1][5] ), .C(\key_mem[2][5] ), 
        .D(\key_mem[3][5] ), .S0(n1404), .S1(n1301), .Y(n102) );
  MXI4X1 U4929 ( .A(n300), .B(n301), .C(n302), .D(n303), .S0(n1271), .S1(n1286), .Y(round_key[37]) );
  MXI4X1 U4930 ( .A(\key_mem[4][37] ), .B(\key_mem[5][37] ), .C(
        \key_mem[6][37] ), .D(\key_mem[7][37] ), .S0(n1357), .S1(n1347), .Y(
        n302) );
  MXI3X1 U4931 ( .A(\key_mem[12][37] ), .B(\key_mem[13][37] ), .C(n297), .S0(
        n1375), .S1(n1340), .Y(n303) );
  MXI4X1 U4932 ( .A(\key_mem[0][37] ), .B(\key_mem[1][37] ), .C(
        \key_mem[2][37] ), .D(\key_mem[3][37] ), .S0(n1359), .S1(n1307), .Y(
        n300) );
  MXI4X1 U4933 ( .A(n460), .B(n461), .C(n462), .D(n463), .S0(n1277), .S1(n1290), .Y(round_key[69]) );
  MXI4X1 U4934 ( .A(\key_mem[4][69] ), .B(\key_mem[5][69] ), .C(
        \key_mem[6][69] ), .D(\key_mem[7][69] ), .S0(n1386), .S1(n1317), .Y(
        n462) );
  MXI3X1 U4935 ( .A(\key_mem[12][69] ), .B(\key_mem[13][69] ), .C(n459), .S0(
        n1374), .S1(n1343), .Y(n463) );
  MXI4X1 U4936 ( .A(\key_mem[0][69] ), .B(\key_mem[1][69] ), .C(
        \key_mem[2][69] ), .D(\key_mem[3][69] ), .S0(n1386), .S1(n1317), .Y(
        n460) );
  MXI4X1 U4937 ( .A(n935), .B(n936), .C(n939), .D(n940), .S0(n1274), .S1(n1280), .Y(round_key[101]) );
  MXI4X1 U4938 ( .A(\key_mem[4][101] ), .B(\key_mem[5][101] ), .C(
        \key_mem[6][101] ), .D(\key_mem[7][101] ), .S0(n1396), .S1(n1327), .Y(
        n939) );
  MXI3X1 U4939 ( .A(\key_mem[12][101] ), .B(\key_mem[13][101] ), .C(n932), 
        .S0(n1374), .S1(n1346), .Y(n940) );
  MXI4X1 U4940 ( .A(\key_mem[0][101] ), .B(\key_mem[1][101] ), .C(
        \key_mem[2][101] ), .D(\key_mem[3][101] ), .S0(n1396), .S1(n1319), .Y(
        n935) );
  MXI4X1 U4941 ( .A(n97), .B(n98), .C(n99), .D(n100), .S0(n1268), .S1(n1283), 
        .Y(round_key[4]) );
  MXI4X1 U4942 ( .A(\key_mem[4][4] ), .B(\key_mem[5][4] ), .C(\key_mem[6][4] ), 
        .D(\key_mem[7][4] ), .S0(n1404), .S1(n1298), .Y(n99) );
  MXI3X1 U4943 ( .A(\key_mem[12][4] ), .B(\key_mem[13][4] ), .C(n96), .S0(
        n1372), .S1(n1337), .Y(n100) );
  MXI4X1 U4944 ( .A(\key_mem[0][4] ), .B(\key_mem[1][4] ), .C(\key_mem[2][4] ), 
        .D(\key_mem[3][4] ), .S0(n1404), .S1(n1299), .Y(n97) );
  MXI4X1 U4945 ( .A(n290), .B(n292), .C(n294), .D(n296), .S0(n1271), .S1(n1286), .Y(round_key[36]) );
  MXI4X1 U4946 ( .A(\key_mem[4][36] ), .B(\key_mem[5][36] ), .C(
        \key_mem[6][36] ), .D(\key_mem[7][36] ), .S0(N31), .S1(n1309), .Y(n294) );
  MXI3X1 U4947 ( .A(\key_mem[12][36] ), .B(\key_mem[13][36] ), .C(n288), .S0(
        n1374), .S1(n1340), .Y(n296) );
  MXI4X1 U4948 ( .A(\key_mem[0][36] ), .B(\key_mem[1][36] ), .C(
        \key_mem[2][36] ), .D(\key_mem[3][36] ), .S0(n1352), .S1(n1309), .Y(
        n290) );
  MXI4X1 U4949 ( .A(n1004), .B(n1007), .C(n1011), .D(n1015), .S0(n1275), .S1(
        N33), .Y(round_key[108]) );
  MXI4X1 U4950 ( .A(\key_mem[4][108] ), .B(\key_mem[5][108] ), .C(
        \key_mem[6][108] ), .D(\key_mem[7][108] ), .S0(n1394), .S1(n1320), .Y(
        n1011) );
  MXI3X1 U4951 ( .A(\key_mem[12][108] ), .B(\key_mem[13][108] ), .C(n1003), 
        .S0(n1376), .S1(n1335), .Y(n1015) );
  MXI4X1 U4952 ( .A(\key_mem[0][108] ), .B(\key_mem[1][108] ), .C(
        \key_mem[2][108] ), .D(\key_mem[3][108] ), .S0(n1394), .S1(n1319), .Y(
        n1004) );
  MXI4X1 U4953 ( .A(n450), .B(n451), .C(n452), .D(n453), .S0(n1265), .S1(n1291), .Y(round_key[67]) );
  MXI4X1 U4954 ( .A(\key_mem[4][67] ), .B(\key_mem[5][67] ), .C(
        \key_mem[6][67] ), .D(\key_mem[7][67] ), .S0(n1387), .S1(n1316), .Y(
        n452) );
  MXI3X1 U4955 ( .A(\key_mem[12][67] ), .B(\key_mem[13][67] ), .C(n449), .S0(
        n1375), .S1(n1343), .Y(n453) );
  MXI4X1 U4956 ( .A(\key_mem[0][67] ), .B(\key_mem[1][67] ), .C(
        \key_mem[2][67] ), .D(\key_mem[3][67] ), .S0(n1387), .S1(n1316), .Y(
        n450) );
  MXI4X1 U4957 ( .A(n330), .B(n331), .C(n332), .D(n333), .S0(n1272), .S1(n1287), .Y(round_key[43]) );
  MXI4X1 U4958 ( .A(\key_mem[4][43] ), .B(\key_mem[5][43] ), .C(
        \key_mem[6][43] ), .D(\key_mem[7][43] ), .S0(n1414), .S1(n1298), .Y(
        n332) );
  MXI3X1 U4959 ( .A(\key_mem[12][43] ), .B(\key_mem[13][43] ), .C(n329), .S0(
        n1379), .S1(n1340), .Y(n333) );
  MXI4X1 U4960 ( .A(\key_mem[0][43] ), .B(\key_mem[1][43] ), .C(
        \key_mem[2][43] ), .D(\key_mem[3][43] ), .S0(n1414), .S1(n1308), .Y(
        n330) );
  MXI4X1 U4961 ( .A(n87), .B(n88), .C(n89), .D(n90), .S0(n1268), .S1(n1283), 
        .Y(round_key[2]) );
  MXI4X1 U4962 ( .A(\key_mem[4][2] ), .B(\key_mem[5][2] ), .C(\key_mem[6][2] ), 
        .D(\key_mem[7][2] ), .S0(n1403), .S1(n1302), .Y(n89) );
  MXI3X1 U4963 ( .A(\key_mem[12][2] ), .B(\key_mem[13][2] ), .C(n86), .S0(
        n1372), .S1(n1336), .Y(n90) );
  MXI4X1 U4964 ( .A(\key_mem[0][2] ), .B(\key_mem[1][2] ), .C(\key_mem[2][2] ), 
        .D(\key_mem[3][2] ), .S0(n1403), .S1(n1308), .Y(n87) );
  MXI4X1 U4965 ( .A(n271), .B(n272), .C(n273), .D(n274), .S0(n1271), .S1(n1286), .Y(round_key[34]) );
  MXI4X1 U4966 ( .A(\key_mem[4][34] ), .B(\key_mem[5][34] ), .C(
        \key_mem[6][34] ), .D(\key_mem[7][34] ), .S0(n1363), .S1(n1309), .Y(
        n273) );
  MXI3X1 U4967 ( .A(\key_mem[12][34] ), .B(\key_mem[13][34] ), .C(n270), .S0(
        n1374), .S1(n1340), .Y(n274) );
  MXI4X1 U4968 ( .A(\key_mem[0][34] ), .B(\key_mem[1][34] ), .C(
        \key_mem[2][34] ), .D(\key_mem[3][34] ), .S0(n1353), .S1(n1331), .Y(
        n271) );
  MXI4X1 U4969 ( .A(n82), .B(n83), .C(n84), .D(n85), .S0(n1265), .S1(n1283), 
        .Y(round_key[1]) );
  MXI4X1 U4970 ( .A(\key_mem[4][1] ), .B(\key_mem[5][1] ), .C(\key_mem[6][1] ), 
        .D(\key_mem[7][1] ), .S0(n1403), .S1(n1295), .Y(n84) );
  MXI3X1 U4971 ( .A(\key_mem[12][1] ), .B(\key_mem[13][1] ), .C(n81), .S0(
        n1372), .S1(n1346), .Y(n85) );
  MXI4X1 U4972 ( .A(\key_mem[0][1] ), .B(\key_mem[1][1] ), .C(\key_mem[2][1] ), 
        .D(\key_mem[3][1] ), .S0(n1403), .S1(n1301), .Y(n82) );
  MXI4X1 U4973 ( .A(n975), .B(n976), .C(n979), .D(n980), .S0(n1274), .S1(n1292), .Y(round_key[105]) );
  MXI4X1 U4974 ( .A(\key_mem[4][105] ), .B(\key_mem[5][105] ), .C(
        \key_mem[6][105] ), .D(\key_mem[7][105] ), .S0(n1395), .S1(n1324), .Y(
        n979) );
  MXI3X1 U4975 ( .A(\key_mem[12][105] ), .B(\key_mem[13][105] ), .C(n972), 
        .S0(n1375), .S1(n1334), .Y(n980) );
  MXI4X1 U4976 ( .A(\key_mem[0][105] ), .B(\key_mem[1][105] ), .C(
        \key_mem[2][105] ), .D(\key_mem[3][105] ), .S0(n1395), .S1(n1324), .Y(
        n975) );
  MXI4X1 U4977 ( .A(n315), .B(n316), .C(n317), .D(n318), .S0(n1272), .S1(n1287), .Y(round_key[40]) );
  MXI4X1 U4978 ( .A(\key_mem[4][40] ), .B(\key_mem[5][40] ), .C(
        \key_mem[6][40] ), .D(\key_mem[7][40] ), .S0(n1415), .S1(n1304), .Y(
        n317) );
  MXI3X1 U4979 ( .A(\key_mem[12][40] ), .B(\key_mem[13][40] ), .C(n314), .S0(
        n1376), .S1(n1340), .Y(n318) );
  MXI4X1 U4980 ( .A(\key_mem[0][40] ), .B(\key_mem[1][40] ), .C(
        \key_mem[2][40] ), .D(\key_mem[3][40] ), .S0(n1415), .S1(n1348), .Y(
        n315) );
  MXI4X1 U4981 ( .A(n964), .B(n967), .C(n968), .D(n971), .S0(n1274), .S1(n1290), .Y(round_key[104]) );
  MXI4X1 U4982 ( .A(\key_mem[4][104] ), .B(\key_mem[5][104] ), .C(
        \key_mem[6][104] ), .D(\key_mem[7][104] ), .S0(n1395), .S1(n1326), .Y(
        n968) );
  MXI3X1 U4983 ( .A(\key_mem[12][104] ), .B(\key_mem[13][104] ), .C(n963), 
        .S0(n1375), .S1(n1335), .Y(n971) );
  MXI4X1 U4984 ( .A(\key_mem[0][104] ), .B(\key_mem[1][104] ), .C(
        \key_mem[2][104] ), .D(\key_mem[3][104] ), .S0(n1395), .S1(n1325), .Y(
        n964) );
  MXI4X1 U4985 ( .A(n261), .B(n262), .C(n263), .D(n264), .S0(n1271), .S1(n1286), .Y(round_key[32]) );
  MXI4X1 U4986 ( .A(\key_mem[4][32] ), .B(\key_mem[5][32] ), .C(
        \key_mem[6][32] ), .D(\key_mem[7][32] ), .S0(n1350), .S1(n1331), .Y(
        n263) );
  MXI3X1 U4987 ( .A(\key_mem[12][32] ), .B(\key_mem[13][32] ), .C(n260), .S0(
        n1373), .S1(n1339), .Y(n264) );
  MXI4X1 U4988 ( .A(\key_mem[0][32] ), .B(\key_mem[1][32] ), .C(
        \key_mem[2][32] ), .D(\key_mem[3][32] ), .S0(n1364), .S1(n1332), .Y(
        n261) );
  MXI4X1 U4989 ( .A(n375), .B(n376), .C(n377), .D(n378), .S0(n1273), .S1(n1288), .Y(round_key[52]) );
  MXI4X1 U4990 ( .A(\key_mem[4][52] ), .B(\key_mem[5][52] ), .C(
        \key_mem[6][52] ), .D(\key_mem[7][52] ), .S0(n1411), .S1(n1310), .Y(
        n377) );
  MXI3X1 U4991 ( .A(\key_mem[12][52] ), .B(\key_mem[13][52] ), .C(n374), .S0(
        n1378), .S1(n1341), .Y(n378) );
  MXI4X1 U4992 ( .A(\key_mem[0][52] ), .B(\key_mem[1][52] ), .C(
        \key_mem[2][52] ), .D(\key_mem[3][52] ), .S0(n1411), .S1(n1311), .Y(
        n375) );
  MXI4X1 U4993 ( .A(n370), .B(n371), .C(n372), .D(n373), .S0(n1273), .S1(n1288), .Y(round_key[51]) );
  MXI4X1 U4994 ( .A(\key_mem[4][51] ), .B(\key_mem[5][51] ), .C(
        \key_mem[6][51] ), .D(\key_mem[7][51] ), .S0(n1411), .S1(n1310), .Y(
        n372) );
  MXI3X1 U4995 ( .A(\key_mem[12][51] ), .B(\key_mem[13][51] ), .C(n369), .S0(
        n1379), .S1(n1341), .Y(n373) );
  MXI4X1 U4996 ( .A(\key_mem[0][51] ), .B(\key_mem[1][51] ), .C(
        \key_mem[2][51] ), .D(\key_mem[3][51] ), .S0(n1411), .S1(n1310), .Y(
        n370) );
  MXI4X1 U4997 ( .A(n365), .B(n366), .C(n367), .D(n368), .S0(n1273), .S1(n1288), .Y(round_key[50]) );
  MXI4X1 U4998 ( .A(\key_mem[4][50] ), .B(\key_mem[5][50] ), .C(
        \key_mem[6][50] ), .D(\key_mem[7][50] ), .S0(n1412), .S1(n1310), .Y(
        n367) );
  MXI3X1 U4999 ( .A(\key_mem[12][50] ), .B(\key_mem[13][50] ), .C(n364), .S0(
        n1378), .S1(n1341), .Y(n368) );
  MXI4X1 U5000 ( .A(\key_mem[0][50] ), .B(\key_mem[1][50] ), .C(
        \key_mem[2][50] ), .D(\key_mem[3][50] ), .S0(n1412), .S1(n1310), .Y(
        n365) );
  MXI4X1 U5001 ( .A(n360), .B(n361), .C(n362), .D(n363), .S0(n1273), .S1(n1288), .Y(round_key[49]) );
  MXI4X1 U5002 ( .A(\key_mem[4][49] ), .B(\key_mem[5][49] ), .C(
        \key_mem[6][49] ), .D(\key_mem[7][49] ), .S0(n1412), .S1(n1309), .Y(
        n362) );
  MXI3X1 U5003 ( .A(\key_mem[12][49] ), .B(\key_mem[13][49] ), .C(n359), .S0(
        n1379), .S1(n1341), .Y(n363) );
  MXI4X1 U5004 ( .A(\key_mem[0][49] ), .B(\key_mem[1][49] ), .C(
        \key_mem[2][49] ), .D(\key_mem[3][49] ), .S0(n1412), .S1(n1309), .Y(
        n360) );
  MXI4X1 U5005 ( .A(n485), .B(n486), .C(n487), .D(n488), .S0(n1269), .S1(n1282), .Y(round_key[74]) );
  MXI4X1 U5006 ( .A(\key_mem[4][74] ), .B(\key_mem[5][74] ), .C(
        \key_mem[6][74] ), .D(\key_mem[7][74] ), .S0(n1384), .S1(n1319), .Y(
        n487) );
  MXI3X1 U5007 ( .A(\key_mem[12][74] ), .B(\key_mem[13][74] ), .C(n484), .S0(
        n1372), .S1(n1344), .Y(n488) );
  MXI4X1 U5008 ( .A(\key_mem[0][74] ), .B(\key_mem[1][74] ), .C(
        \key_mem[2][74] ), .D(\key_mem[3][74] ), .S0(n1384), .S1(n1319), .Y(
        n485) );
  MXI4X1 U5009 ( .A(n480), .B(n481), .C(n482), .D(n483), .S0(n1267), .S1(n1292), .Y(round_key[73]) );
  MXI4X1 U5010 ( .A(\key_mem[4][73] ), .B(\key_mem[5][73] ), .C(
        \key_mem[6][73] ), .D(\key_mem[7][73] ), .S0(n1384), .S1(n1318), .Y(
        n482) );
  MXI3X1 U5011 ( .A(\key_mem[12][73] ), .B(\key_mem[13][73] ), .C(n479), .S0(
        n1372), .S1(n1344), .Y(n483) );
  MXI4X1 U5012 ( .A(\key_mem[0][73] ), .B(\key_mem[1][73] ), .C(
        \key_mem[2][73] ), .D(\key_mem[3][73] ), .S0(n1384), .S1(n1318), .Y(
        n480) );
  MXI4X1 U5013 ( .A(n924), .B(n927), .C(n928), .D(n931), .S0(n1274), .S1(n1290), .Y(round_key[100]) );
  MXI4X1 U5014 ( .A(\key_mem[4][100] ), .B(\key_mem[5][100] ), .C(
        \key_mem[6][100] ), .D(\key_mem[7][100] ), .S0(n1396), .S1(n1327), .Y(
        n928) );
  MXI3X1 U5015 ( .A(\key_mem[12][100] ), .B(\key_mem[13][100] ), .C(n923), 
        .S0(n1374), .S1(n1346), .Y(n931) );
  MXI4X1 U5016 ( .A(\key_mem[0][100] ), .B(\key_mem[1][100] ), .C(
        \key_mem[2][100] ), .D(\key_mem[3][100] ), .S0(n1396), .S1(n1327), .Y(
        n924) );
  MXI4X1 U5017 ( .A(n915), .B(n916), .C(n919), .D(n920), .S0(n1274), .S1(n1283), .Y(round_key[99]) );
  MXI4X1 U5018 ( .A(\key_mem[4][99] ), .B(\key_mem[5][99] ), .C(
        \key_mem[6][99] ), .D(\key_mem[7][99] ), .S0(n1397), .S1(N32), .Y(n919) );
  MXI3X1 U5019 ( .A(\key_mem[12][99] ), .B(\key_mem[13][99] ), .C(n912), .S0(
        n1374), .S1(n1346), .Y(n920) );
  MXI4X1 U5020 ( .A(\key_mem[0][99] ), .B(\key_mem[1][99] ), .C(
        \key_mem[2][99] ), .D(\key_mem[3][99] ), .S0(n1396), .S1(N32), .Y(n915) );
  MXI4X1 U5021 ( .A(n876), .B(n907), .C(n908), .D(n911), .S0(n1274), .S1(n1280), .Y(round_key[98]) );
  MXI4X1 U5022 ( .A(\key_mem[4][98] ), .B(\key_mem[5][98] ), .C(
        \key_mem[6][98] ), .D(\key_mem[7][98] ), .S0(n1397), .S1(n1348), .Y(
        n908) );
  MXI3X1 U5023 ( .A(\key_mem[12][98] ), .B(\key_mem[13][98] ), .C(n875), .S0(
        n1373), .S1(n1346), .Y(n911) );
  MXI4X1 U5024 ( .A(\key_mem[0][98] ), .B(\key_mem[1][98] ), .C(
        \key_mem[2][98] ), .D(\key_mem[3][98] ), .S0(n1397), .S1(n1347), .Y(
        n876) );
  MXI4X1 U5025 ( .A(n747), .B(n748), .C(n751), .D(n755), .S0(n1266), .S1(n1280), .Y(round_key[96]) );
  MXI4X1 U5026 ( .A(\key_mem[4][96] ), .B(\key_mem[5][96] ), .C(
        \key_mem[6][96] ), .D(\key_mem[7][96] ), .S0(n1397), .S1(N32), .Y(n751) );
  MXI3X1 U5027 ( .A(\key_mem[12][96] ), .B(\key_mem[13][96] ), .C(n746), .S0(
        n1373), .S1(n1346), .Y(n755) );
  MXI4X1 U5028 ( .A(\key_mem[0][96] ), .B(\key_mem[1][96] ), .C(
        \key_mem[2][96] ), .D(\key_mem[3][96] ), .S0(n1397), .S1(n1347), .Y(
        n747) );
  MXI4X1 U5029 ( .A(n550), .B(n551), .C(n552), .D(n553), .S0(n1269), .S1(n1291), .Y(round_key[87]) );
  MXI3X1 U5030 ( .A(\key_mem[12][87] ), .B(\key_mem[13][87] ), .C(n549), .S0(
        n1370), .S1(n1345), .Y(n553) );
  MXI4X1 U5031 ( .A(\key_mem[4][87] ), .B(\key_mem[5][87] ), .C(
        \key_mem[6][87] ), .D(\key_mem[7][87] ), .S0(n1400), .S1(n1324), .Y(
        n552) );
  MXI4X1 U5032 ( .A(\key_mem[0][87] ), .B(\key_mem[1][87] ), .C(
        \key_mem[2][87] ), .D(\key_mem[3][87] ), .S0(n1400), .S1(n1324), .Y(
        n550) );
  MXI4X1 U5033 ( .A(n390), .B(n391), .C(n392), .D(n393), .S0(n1273), .S1(n1288), .Y(round_key[55]) );
  MXI4X1 U5034 ( .A(\key_mem[4][55] ), .B(\key_mem[5][55] ), .C(
        \key_mem[6][55] ), .D(\key_mem[7][55] ), .S0(n1380), .S1(n1312), .Y(
        n392) );
  MXI3X1 U5035 ( .A(\key_mem[12][55] ), .B(\key_mem[13][55] ), .C(n389), .S0(
        n1376), .S1(n1342), .Y(n393) );
  MXI4X1 U5036 ( .A(\key_mem[0][55] ), .B(\key_mem[1][55] ), .C(
        \key_mem[2][55] ), .D(\key_mem[3][55] ), .S0(n1381), .S1(n1312), .Y(
        n390) );
  MXI4X1 U5037 ( .A(n206), .B(n207), .C(n208), .D(n209), .S0(n1270), .S1(n1285), .Y(round_key[21]) );
  MXI3X1 U5038 ( .A(\key_mem[12][21] ), .B(\key_mem[13][21] ), .C(n205), .S0(
        n1369), .S1(n1338), .Y(n209) );
  MXI4X1 U5039 ( .A(\key_mem[4][21] ), .B(\key_mem[5][21] ), .C(
        \key_mem[6][21] ), .D(\key_mem[7][21] ), .S0(n1409), .S1(n1308), .Y(
        n208) );
  MXI4X1 U5040 ( .A(\key_mem[0][21] ), .B(\key_mem[1][21] ), .C(
        \key_mem[2][21] ), .D(\key_mem[3][21] ), .S0(n1409), .S1(n1307), .Y(
        n206) );
  MXI4X1 U5041 ( .A(n201), .B(n202), .C(n203), .D(n204), .S0(n1270), .S1(n1285), .Y(round_key[20]) );
  MXI3X1 U5042 ( .A(\key_mem[12][20] ), .B(\key_mem[13][20] ), .C(n200), .S0(
        n1369), .S1(n1338), .Y(n204) );
  MXI4X1 U5043 ( .A(\key_mem[4][20] ), .B(\key_mem[5][20] ), .C(
        \key_mem[6][20] ), .D(\key_mem[7][20] ), .S0(n1408), .S1(n1296), .Y(
        n203) );
  MXI4X1 U5044 ( .A(\key_mem[0][20] ), .B(\key_mem[1][20] ), .C(
        \key_mem[2][20] ), .D(\key_mem[3][20] ), .S0(n1408), .S1(n1293), .Y(
        n201) );
  MXI4X1 U5045 ( .A(n530), .B(n531), .C(n532), .D(n533), .S0(n1267), .S1(n1291), .Y(round_key[83]) );
  MXI3X1 U5046 ( .A(\key_mem[12][83] ), .B(\key_mem[13][83] ), .C(n529), .S0(
        n1369), .S1(n1345), .Y(n533) );
  MXI4X1 U5047 ( .A(\key_mem[4][83] ), .B(\key_mem[5][83] ), .C(
        \key_mem[6][83] ), .D(\key_mem[7][83] ), .S0(n1401), .S1(n1322), .Y(
        n532) );
  MXI4X1 U5048 ( .A(\key_mem[0][83] ), .B(\key_mem[1][83] ), .C(
        \key_mem[2][83] ), .D(\key_mem[3][83] ), .S0(n1401), .S1(n1322), .Y(
        n530) );
  MXI4X1 U5049 ( .A(n545), .B(n546), .C(n547), .D(n548), .S0(n1278), .S1(n1282), .Y(round_key[86]) );
  MXI3X1 U5050 ( .A(\key_mem[12][86] ), .B(\key_mem[13][86] ), .C(n544), .S0(
        n1357), .S1(n1345), .Y(n548) );
  MXI4X1 U5051 ( .A(\key_mem[4][86] ), .B(\key_mem[5][86] ), .C(
        \key_mem[6][86] ), .D(\key_mem[7][86] ), .S0(n1400), .S1(n1323), .Y(
        n547) );
  MXI4X1 U5052 ( .A(\key_mem[0][86] ), .B(\key_mem[1][86] ), .C(
        \key_mem[2][86] ), .D(\key_mem[3][86] ), .S0(n1400), .S1(n1323), .Y(
        n545) );
  MXI4X1 U5053 ( .A(n127), .B(n128), .C(n129), .D(n130), .S0(n1268), .S1(n1284), .Y(round_key[10]) );
  MXI3X1 U5054 ( .A(\key_mem[12][10] ), .B(\key_mem[13][10] ), .C(n126), .S0(
        n1370), .S1(n1337), .Y(n130) );
  MXI4X1 U5055 ( .A(\key_mem[4][10] ), .B(\key_mem[5][10] ), .C(
        \key_mem[6][10] ), .D(\key_mem[7][10] ), .S0(n1405), .S1(n1328), .Y(
        n129) );
  MXI4X1 U5056 ( .A(\key_mem[0][10] ), .B(\key_mem[1][10] ), .C(
        \key_mem[2][10] ), .D(\key_mem[3][10] ), .S0(n1405), .S1(n1328), .Y(
        n127) );
  MXI4X1 U5057 ( .A(n122), .B(n123), .C(n124), .D(n125), .S0(n1278), .S1(n1284), .Y(round_key[9]) );
  MXI3X1 U5058 ( .A(\key_mem[12][9] ), .B(\key_mem[13][9] ), .C(n121), .S0(
        n1370), .S1(n1337), .Y(n125) );
  MXI4X1 U5059 ( .A(\key_mem[4][9] ), .B(\key_mem[5][9] ), .C(\key_mem[6][9] ), 
        .D(\key_mem[7][9] ), .S0(n1405), .S1(n1328), .Y(n124) );
  MXI4X1 U5060 ( .A(\key_mem[0][9] ), .B(\key_mem[1][9] ), .C(\key_mem[2][9] ), 
        .D(\key_mem[3][9] ), .S0(n1405), .S1(n1328), .Y(n122) );
  MXI4X1 U5061 ( .A(n107), .B(n108), .C(n109), .D(n110), .S0(n1266), .S1(n1283), .Y(round_key[6]) );
  MXI4X1 U5062 ( .A(\key_mem[4][6] ), .B(\key_mem[5][6] ), .C(\key_mem[6][6] ), 
        .D(\key_mem[7][6] ), .S0(n1404), .S1(n1304), .Y(n109) );
  MXI3X1 U5063 ( .A(\key_mem[12][6] ), .B(\key_mem[13][6] ), .C(n106), .S0(
        n1371), .S1(n1337), .Y(n110) );
  MXI4X1 U5064 ( .A(\key_mem[0][6] ), .B(\key_mem[1][6] ), .C(\key_mem[2][6] ), 
        .D(\key_mem[3][6] ), .S0(n1404), .S1(n1296), .Y(n107) );
  MXI4X1 U5065 ( .A(n455), .B(n456), .C(n457), .D(n458), .S0(n1266), .S1(n1279), .Y(round_key[68]) );
  MXI4X1 U5066 ( .A(\key_mem[4][68] ), .B(\key_mem[5][68] ), .C(
        \key_mem[6][68] ), .D(\key_mem[7][68] ), .S0(n1387), .S1(n1316), .Y(
        n457) );
  MXI3X1 U5067 ( .A(\key_mem[12][68] ), .B(\key_mem[13][68] ), .C(n454), .S0(
        n1375), .S1(n1343), .Y(n458) );
  MXI4X1 U5068 ( .A(\key_mem[0][68] ), .B(\key_mem[1][68] ), .C(
        \key_mem[2][68] ), .D(\key_mem[3][68] ), .S0(n1387), .S1(n1317), .Y(
        n455) );
  MXI4X1 U5069 ( .A(n335), .B(n336), .C(n337), .D(n338), .S0(n1272), .S1(n1287), .Y(round_key[44]) );
  MXI4X1 U5070 ( .A(\key_mem[4][44] ), .B(\key_mem[5][44] ), .C(
        \key_mem[6][44] ), .D(\key_mem[7][44] ), .S0(n1413), .S1(n1302), .Y(
        n337) );
  MXI3X1 U5071 ( .A(\key_mem[12][44] ), .B(\key_mem[13][44] ), .C(n334), .S0(
        n1379), .S1(n1341), .Y(n338) );
  MXI4X1 U5072 ( .A(\key_mem[0][44] ), .B(\key_mem[1][44] ), .C(
        \key_mem[2][44] ), .D(\key_mem[3][44] ), .S0(n1413), .S1(n1305), .Y(
        n335) );
  MXI4X1 U5073 ( .A(n92), .B(n93), .C(n94), .D(n95), .S0(n1278), .S1(n1283), 
        .Y(round_key[3]) );
  MXI4X1 U5074 ( .A(\key_mem[4][3] ), .B(\key_mem[5][3] ), .C(\key_mem[6][3] ), 
        .D(\key_mem[7][3] ), .S0(n1403), .S1(n1293), .Y(n94) );
  MXI3X1 U5075 ( .A(\key_mem[12][3] ), .B(\key_mem[13][3] ), .C(n91), .S0(
        n1372), .S1(n1336), .Y(n95) );
  MXI4X1 U5076 ( .A(\key_mem[0][3] ), .B(\key_mem[1][3] ), .C(\key_mem[2][3] ), 
        .D(\key_mem[3][3] ), .S0(n1403), .S1(n1308), .Y(n92) );
  MXI4X1 U5077 ( .A(n325), .B(n326), .C(n327), .D(n328), .S0(n1272), .S1(n1287), .Y(round_key[42]) );
  MXI4X1 U5078 ( .A(\key_mem[4][42] ), .B(\key_mem[5][42] ), .C(
        \key_mem[6][42] ), .D(\key_mem[7][42] ), .S0(n1414), .S1(n1302), .Y(
        n327) );
  MXI3X1 U5079 ( .A(\key_mem[12][42] ), .B(\key_mem[13][42] ), .C(n324), .S0(
        n1377), .S1(n1340), .Y(n328) );
  MXI4X1 U5080 ( .A(\key_mem[0][42] ), .B(\key_mem[1][42] ), .C(
        \key_mem[2][42] ), .D(\key_mem[3][42] ), .S0(n1414), .S1(n1298), .Y(
        n325) );
  MXI4X1 U5081 ( .A(n984), .B(n987), .C(n988), .D(n991), .S0(n1274), .S1(n1290), .Y(round_key[106]) );
  MXI4X1 U5082 ( .A(\key_mem[4][106] ), .B(\key_mem[5][106] ), .C(
        \key_mem[6][106] ), .D(\key_mem[7][106] ), .S0(n1394), .S1(n1323), .Y(
        n988) );
  MXI3X1 U5083 ( .A(\key_mem[12][106] ), .B(\key_mem[13][106] ), .C(n983), 
        .S0(n1375), .S1(n1334), .Y(n991) );
  MXI4X1 U5084 ( .A(\key_mem[0][106] ), .B(\key_mem[1][106] ), .C(
        \key_mem[2][106] ), .D(\key_mem[3][106] ), .S0(n1394), .S1(n1322), .Y(
        n984) );
  MXI4X1 U5085 ( .A(n445), .B(n446), .C(n447), .D(n448), .S0(n1266), .S1(n1280), .Y(round_key[66]) );
  MXI4X1 U5086 ( .A(\key_mem[4][66] ), .B(\key_mem[5][66] ), .C(
        \key_mem[6][66] ), .D(\key_mem[7][66] ), .S0(n1388), .S1(n1316), .Y(
        n447) );
  MXI3X1 U5087 ( .A(\key_mem[12][66] ), .B(\key_mem[13][66] ), .C(n444), .S0(
        n1377), .S1(n1343), .Y(n448) );
  MXI4X1 U5088 ( .A(\key_mem[0][66] ), .B(\key_mem[1][66] ), .C(
        \key_mem[2][66] ), .D(\key_mem[3][66] ), .S0(n1388), .S1(n1316), .Y(
        n445) );
  MXI4X1 U5089 ( .A(n266), .B(n267), .C(n268), .D(n269), .S0(n1271), .S1(n1286), .Y(round_key[33]) );
  MXI4X1 U5090 ( .A(\key_mem[4][33] ), .B(\key_mem[5][33] ), .C(
        \key_mem[6][33] ), .D(\key_mem[7][33] ), .S0(n1417), .S1(n1331), .Y(
        n268) );
  MXI3X1 U5091 ( .A(\key_mem[12][33] ), .B(\key_mem[13][33] ), .C(n265), .S0(
        n1374), .S1(n1339), .Y(n269) );
  MXI4X1 U5092 ( .A(\key_mem[0][33] ), .B(\key_mem[1][33] ), .C(
        \key_mem[2][33] ), .D(\key_mem[3][33] ), .S0(n1351), .S1(n1331), .Y(
        n266) );
  MXI4X1 U5093 ( .A(n440), .B(n441), .C(n442), .D(n443), .S0(n1265), .S1(n1292), .Y(round_key[65]) );
  MXI4X1 U5094 ( .A(\key_mem[4][65] ), .B(\key_mem[5][65] ), .C(
        \key_mem[6][65] ), .D(\key_mem[7][65] ), .S0(n1388), .S1(n1315), .Y(
        n442) );
  MXI3X1 U5095 ( .A(\key_mem[12][65] ), .B(\key_mem[13][65] ), .C(n439), .S0(
        n1377), .S1(n1343), .Y(n443) );
  MXI4X1 U5096 ( .A(\key_mem[0][65] ), .B(\key_mem[1][65] ), .C(
        \key_mem[2][65] ), .D(\key_mem[3][65] ), .S0(n1388), .S1(n1315), .Y(
        n440) );
  MXI4X1 U5097 ( .A(n320), .B(n321), .C(n322), .D(n323), .S0(n1272), .S1(n1287), .Y(round_key[41]) );
  MXI4X1 U5098 ( .A(\key_mem[4][41] ), .B(\key_mem[5][41] ), .C(
        \key_mem[6][41] ), .D(\key_mem[7][41] ), .S0(n1414), .S1(n1297), .Y(
        n322) );
  MXI3X1 U5099 ( .A(\key_mem[12][41] ), .B(\key_mem[13][41] ), .C(n319), .S0(
        n1376), .S1(n1340), .Y(n323) );
  MXI4X1 U5100 ( .A(\key_mem[0][41] ), .B(\key_mem[1][41] ), .C(
        \key_mem[2][41] ), .D(\key_mem[3][41] ), .S0(n1414), .S1(n1297), .Y(
        n320) );
  MXI4X1 U5101 ( .A(n77), .B(n78), .C(n79), .D(n80), .S0(n1266), .S1(n1283), 
        .Y(round_key[0]) );
  MXI4X1 U5102 ( .A(\key_mem[4][0] ), .B(\key_mem[5][0] ), .C(\key_mem[6][0] ), 
        .D(\key_mem[7][0] ), .S0(n1402), .S1(n1327), .Y(n79) );
  MXI3X1 U5103 ( .A(\key_mem[12][0] ), .B(\key_mem[13][0] ), .C(n76), .S0(
        n1373), .S1(n1343), .Y(n80) );
  MXI4X1 U5104 ( .A(\key_mem[0][0] ), .B(\key_mem[1][0] ), .C(\key_mem[2][0] ), 
        .D(\key_mem[3][0] ), .S0(n1402), .S1(n1327), .Y(n77) );
  MXI4X1 U5105 ( .A(n355), .B(n356), .C(n357), .D(n358), .S0(n1273), .S1(n1288), .Y(round_key[48]) );
  MXI4X1 U5106 ( .A(n495), .B(n496), .C(n497), .D(n498), .S0(n1278), .S1(n1282), .Y(round_key[76]) );
  MXI3X1 U5107 ( .A(\key_mem[12][76] ), .B(\key_mem[13][76] ), .C(n494), .S0(
        n1370), .S1(n1344), .Y(n498) );
  MXI4X1 U5108 ( .A(\key_mem[4][76] ), .B(\key_mem[5][76] ), .C(
        \key_mem[6][76] ), .D(\key_mem[7][76] ), .S0(n1382), .S1(n1320), .Y(
        n497) );
  MXI4X1 U5109 ( .A(\key_mem[0][76] ), .B(\key_mem[1][76] ), .C(
        \key_mem[2][76] ), .D(\key_mem[3][76] ), .S0(n1382), .S1(n1320), .Y(
        n495) );
  MXI4X1 U5110 ( .A(n763), .B(n767), .C(n771), .D(n775), .S0(n1267), .S1(n1282), .Y(round_key[97]) );
  MXI4X1 U5111 ( .A(\key_mem[4][97] ), .B(\key_mem[5][97] ), .C(
        \key_mem[6][97] ), .D(\key_mem[7][97] ), .S0(n1397), .S1(N32), .Y(n771) );
  MXI3X1 U5112 ( .A(\key_mem[12][97] ), .B(\key_mem[13][97] ), .C(n759), .S0(
        n1373), .S1(n1346), .Y(n775) );
  MXI4X1 U5113 ( .A(\key_mem[0][97] ), .B(\key_mem[1][97] ), .C(
        \key_mem[2][97] ), .D(\key_mem[3][97] ), .S0(n1397), .S1(N32), .Y(n763) );
  MXI4X1 U5114 ( .A(n435), .B(n436), .C(n437), .D(n438), .S0(n1268), .S1(n1283), .Y(round_key[64]) );
  MXI4X1 U5115 ( .A(\key_mem[4][64] ), .B(\key_mem[5][64] ), .C(
        \key_mem[6][64] ), .D(\key_mem[7][64] ), .S0(n1387), .S1(n1315), .Y(
        n437) );
  MXI3X1 U5116 ( .A(\key_mem[12][64] ), .B(\key_mem[13][64] ), .C(n434), .S0(
        n1377), .S1(n1336), .Y(n438) );
  MXI4X1 U5117 ( .A(\key_mem[0][64] ), .B(\key_mem[1][64] ), .C(
        \key_mem[2][64] ), .D(\key_mem[3][64] ), .S0(n1387), .S1(n1315), .Y(
        n435) );
  NOR2BX1 U5118 ( .AN(\key_mem[14][119] ), .B(n1368), .Y(n1187) );
  NOR2BX1 U5119 ( .AN(\key_mem[14][87] ), .B(n1359), .Y(n549) );
  NOR2BX1 U5120 ( .AN(\key_mem[14][55] ), .B(n1357), .Y(n389) );
  NOR2BX1 U5121 ( .AN(\key_mem[14][21] ), .B(n1361), .Y(n205) );
  NOR2BX1 U5122 ( .AN(\key_mem[14][116] ), .B(n1350), .Y(n1151) );
  NOR2BX1 U5123 ( .AN(\key_mem[14][84] ), .B(n1364), .Y(n534) );
  NOR2BX1 U5124 ( .AN(\key_mem[14][20] ), .B(N31), .Y(n200) );
  NOR2BX1 U5125 ( .AN(\key_mem[14][115] ), .B(n1366), .Y(n1132) );
  NOR2BX1 U5126 ( .AN(\key_mem[14][114] ), .B(n1364), .Y(n1120) );
  NOR2BX1 U5127 ( .AN(\key_mem[14][82] ), .B(n1418), .Y(n524) );
  NOR2BX1 U5128 ( .AN(\key_mem[14][18] ), .B(n1351), .Y(n166) );
  NOR2BX1 U5129 ( .AN(\key_mem[14][81] ), .B(n1350), .Y(n519) );
  NOR2BX1 U5130 ( .AN(\key_mem[14][17] ), .B(n1363), .Y(n161) );
  NOR2BX1 U5131 ( .AN(\key_mem[14][113] ), .B(n1358), .Y(n1100) );
  NOR2BX1 U5132 ( .AN(\key_mem[14][80] ), .B(n1365), .Y(n514) );
  NOR2BX1 U5133 ( .AN(\key_mem[14][23] ), .B(n1356), .Y(n215) );
  NOR2BX1 U5134 ( .AN(\key_mem[14][118] ), .B(n1350), .Y(n1176) );
  NOR2BX1 U5135 ( .AN(\key_mem[14][85] ), .B(n1356), .Y(n539) );
  NOR2BX1 U5136 ( .AN(\key_mem[14][53] ), .B(n1359), .Y(n379) );
  NOR2BX1 U5137 ( .AN(\key_mem[14][16] ), .B(n1358), .Y(n156) );
  NOR2BX1 U5138 ( .AN(\key_mem[14][117] ), .B(n1366), .Y(n1167) );
  NOR2BX1 U5139 ( .AN(\key_mem[14][45] ), .B(n1364), .Y(n339) );
  NOR2BX1 U5140 ( .AN(\key_mem[14][109] ), .B(n1358), .Y(n1019) );
  NOR2BX1 U5141 ( .AN(\key_mem[14][86] ), .B(n1352), .Y(n544) );
  NOR2BX1 U5142 ( .AN(\key_mem[14][54] ), .B(n1355), .Y(n384) );
  NOR2BX1 U5143 ( .AN(\key_mem[14][110] ), .B(n1417), .Y(n1040) );
  NOR2BX1 U5144 ( .AN(\key_mem[14][46] ), .B(n1363), .Y(n344) );
  NOR2BX1 U5145 ( .AN(\key_mem[14][22] ), .B(n1362), .Y(n210) );
  NOR2BX1 U5146 ( .AN(\key_mem[14][78] ), .B(n1417), .Y(n504) );
  NOR2BX1 U5147 ( .AN(\key_mem[14][14] ), .B(n1368), .Y(n146) );
  NOR2BX1 U5148 ( .AN(\key_mem[14][77] ), .B(n1359), .Y(n499) );
  NOR2BX1 U5149 ( .AN(\key_mem[14][13] ), .B(n1417), .Y(n141) );
  NOR2BX1 U5150 ( .AN(\key_mem[14][12] ), .B(n1355), .Y(n136) );
  NOR2BX1 U5151 ( .AN(\key_mem[14][10] ), .B(n1366), .Y(n126) );
  NOR2BX1 U5152 ( .AN(\key_mem[14][9] ), .B(n1349), .Y(n121) );
  NOR2BX1 U5153 ( .AN(\key_mem[14][72] ), .B(n1354), .Y(n474) );
  NOR2BX1 U5154 ( .AN(\key_mem[14][8] ), .B(n1361), .Y(n116) );
  NOR2BX1 U5155 ( .AN(\key_mem[14][112] ), .B(n1418), .Y(n1080) );
  NOR2BX1 U5156 ( .AN(\key_mem[14][47] ), .B(n1361), .Y(n349) );
  NOR2BX1 U5157 ( .AN(\key_mem[14][71] ), .B(n1351), .Y(n469) );
  NOR2BX1 U5158 ( .AN(\key_mem[14][15] ), .B(n1367), .Y(n151) );
  NOR2BX1 U5159 ( .AN(\key_mem[14][39] ), .B(n1417), .Y(n309) );
  NOR2BX1 U5160 ( .AN(\key_mem[14][111] ), .B(n1356), .Y(n1060) );
  NOR2BX1 U5161 ( .AN(\key_mem[14][7] ), .B(n1364), .Y(n111) );
  NOR2BX1 U5162 ( .AN(\key_mem[14][79] ), .B(n1357), .Y(n509) );
  NOR2BX1 U5163 ( .AN(\key_mem[14][103] ), .B(n1367), .Y(n952) );
  NOR2BX1 U5164 ( .AN(\key_mem[14][6] ), .B(N31), .Y(n106) );
  NOR2BX1 U5165 ( .AN(\key_mem[14][38] ), .B(n1364), .Y(n304) );
  NOR2BX1 U5166 ( .AN(\key_mem[14][70] ), .B(n1418), .Y(n464) );
  NOR2BX1 U5167 ( .AN(\key_mem[14][102] ), .B(n1367), .Y(n943) );
  NOR2BX1 U5168 ( .AN(\key_mem[14][5] ), .B(n1360), .Y(n101) );
  NOR2BX1 U5169 ( .AN(\key_mem[14][37] ), .B(n1362), .Y(n297) );
  NOR2BX1 U5170 ( .AN(\key_mem[14][69] ), .B(n1354), .Y(n459) );
  NOR2BX1 U5171 ( .AN(\key_mem[14][101] ), .B(n1363), .Y(n932) );
  NOR2BX1 U5172 ( .AN(\key_mem[14][4] ), .B(n1354), .Y(n96) );
  NOR2BX1 U5173 ( .AN(\key_mem[14][36] ), .B(n1354), .Y(n288) );
  NOR2BX1 U5174 ( .AN(\key_mem[14][68] ), .B(n1355), .Y(n454) );
  NOR2BX1 U5175 ( .AN(\key_mem[14][44] ), .B(n1365), .Y(n334) );
  NOR2BX1 U5176 ( .AN(\key_mem[14][108] ), .B(n1368), .Y(n1003) );
  NOR2BX1 U5177 ( .AN(\key_mem[14][42] ), .B(n1360), .Y(n324) );
  NOR2BX1 U5178 ( .AN(\key_mem[14][106] ), .B(n1366), .Y(n983) );
  NOR2BX1 U5179 ( .AN(\key_mem[14][2] ), .B(n1359), .Y(n86) );
  NOR2BX1 U5180 ( .AN(\key_mem[14][34] ), .B(n1416), .Y(n270) );
  NOR2BX1 U5181 ( .AN(\key_mem[14][66] ), .B(n1349), .Y(n444) );
  NOR2BX1 U5182 ( .AN(\key_mem[14][1] ), .B(n1362), .Y(n81) );
  NOR2BX1 U5183 ( .AN(\key_mem[14][33] ), .B(n1416), .Y(n265) );
  NOR2BX1 U5184 ( .AN(\key_mem[14][65] ), .B(n1361), .Y(n439) );
  NOR2BX1 U5185 ( .AN(\key_mem[14][41] ), .B(n1355), .Y(n319) );
  NOR2BX1 U5186 ( .AN(\key_mem[14][105] ), .B(n1351), .Y(n972) );
  NOR2BX1 U5187 ( .AN(\key_mem[14][40] ), .B(n1354), .Y(n314) );
  NOR2BX1 U5188 ( .AN(\key_mem[14][104] ), .B(n1418), .Y(n963) );
  NOR2BX1 U5189 ( .AN(\key_mem[14][0] ), .B(n1416), .Y(n76) );
  NOR2BX1 U5190 ( .AN(\key_mem[14][32] ), .B(n1416), .Y(n260) );
  NOR2BX1 U5191 ( .AN(\key_mem[14][62] ), .B(n1363), .Y(n424) );
  NOR2BX1 U5192 ( .AN(\key_mem[14][29] ), .B(n1416), .Y(n245) );
  NOR2BX1 U5193 ( .AN(\key_mem[14][52] ), .B(n1354), .Y(n374) );
  NOR2BX1 U5194 ( .AN(\key_mem[14][28] ), .B(n1416), .Y(n240) );
  NOR2BX1 U5195 ( .AN(\key_mem[14][27] ), .B(n1416), .Y(n235) );
  NOR2BX1 U5196 ( .AN(\key_mem[14][50] ), .B(n1417), .Y(n364) );
  NOR2BX1 U5197 ( .AN(\key_mem[14][26] ), .B(n1360), .Y(n230) );
  NOR2BX1 U5198 ( .AN(\key_mem[14][49] ), .B(n1361), .Y(n359) );
  NOR2BX1 U5199 ( .AN(\key_mem[14][25] ), .B(n1365), .Y(n225) );
  NOR2BX1 U5200 ( .AN(\key_mem[14][56] ), .B(n1360), .Y(n394) );
  NOR2BX1 U5201 ( .AN(\key_mem[14][61] ), .B(N31), .Y(n419) );
  NOR2BX1 U5202 ( .AN(\key_mem[14][60] ), .B(n1359), .Y(n414) );
  NOR2BX1 U5203 ( .AN(\key_mem[14][59] ), .B(n1361), .Y(n409) );
  NOR2BX1 U5204 ( .AN(\key_mem[14][58] ), .B(n1365), .Y(n404) );
  NOR2BX1 U5205 ( .AN(\key_mem[14][57] ), .B(n1355), .Y(n399) );
  NOR2BX1 U5206 ( .AN(\key_mem[14][24] ), .B(n1363), .Y(n220) );
  NOR2BX1 U5207 ( .AN(\key_mem[14][31] ), .B(n1416), .Y(n255) );
  NOR2BX1 U5208 ( .AN(\key_mem[14][30] ), .B(n1416), .Y(n250) );
  NOR2BX1 U5209 ( .AN(\key_mem[14][126] ), .B(n1367), .Y(n1255) );
  NOR2BX1 U5210 ( .AN(\key_mem[14][125] ), .B(n1350), .Y(n1247) );
  NOR2BX1 U5211 ( .AN(\key_mem[14][124] ), .B(n1349), .Y(n1236) );
  NOR2BX1 U5212 ( .AN(\key_mem[14][122] ), .B(n1366), .Y(n1216) );
  NOR2BX1 U5213 ( .AN(\key_mem[14][121] ), .B(n1367), .Y(n1207) );
  NOR2BX1 U5214 ( .AN(\key_mem[14][120] ), .B(n1358), .Y(n1196) );
  NOR2BX1 U5215 ( .AN(\key_mem[14][127] ), .B(n1360), .Y(n1260) );
  NOR2BX1 U5216 ( .AN(\key_mem[14][94] ), .B(n1417), .Y(n584) );
  NOR2BX1 U5217 ( .AN(\key_mem[14][93] ), .B(n1362), .Y(n579) );
  NOR2BX1 U5218 ( .AN(\key_mem[14][92] ), .B(n1366), .Y(n574) );
  NOR2BX1 U5219 ( .AN(\key_mem[14][91] ), .B(n1357), .Y(n569) );
  NOR2BX1 U5220 ( .AN(\key_mem[14][90] ), .B(n1367), .Y(n564) );
  NOR2BX1 U5221 ( .AN(\key_mem[14][89] ), .B(n1418), .Y(n559) );
  NOR2BX1 U5222 ( .AN(\key_mem[14][88] ), .B(n1358), .Y(n554) );
  NOR2BX1 U5223 ( .AN(\key_mem[14][95] ), .B(n1368), .Y(n589) );
  NOR2BX1 U5224 ( .AN(\key_mem[14][63] ), .B(n1365), .Y(n429) );
  NOR2BX1 U5225 ( .AN(\key_mem[14][76] ), .B(n1368), .Y(n494) );
  NOR2BX1 U5226 ( .AN(\key_mem[14][74] ), .B(n1358), .Y(n484) );
  NOR2BX1 U5227 ( .AN(\key_mem[14][73] ), .B(n1418), .Y(n479) );
  NOR2BX1 U5228 ( .AN(\key_mem[14][100] ), .B(n1357), .Y(n923) );
  NOR2BX1 U5229 ( .AN(\key_mem[14][98] ), .B(n1367), .Y(n875) );
  NOR2BX1 U5230 ( .AN(\key_mem[14][97] ), .B(n1368), .Y(n759) );
  NOR2BX1 U5231 ( .AN(\key_mem[14][64] ), .B(n1355), .Y(n434) );
  NOR2BX1 U5232 ( .AN(\key_mem[14][96] ), .B(n1354), .Y(n746) );
  MXI4X1 U5233 ( .A(\key_mem[8][119] ), .B(\key_mem[9][119] ), .C(
        \key_mem[10][119] ), .D(\key_mem[11][119] ), .S0(n1391), .S1(n1331), 
        .Y(n1191) );
  MXI4X1 U5234 ( .A(\key_mem[8][87] ), .B(\key_mem[9][87] ), .C(
        \key_mem[10][87] ), .D(\key_mem[11][87] ), .S0(n1400), .S1(n1324), .Y(
        n551) );
  MXI4X1 U5235 ( .A(\key_mem[8][55] ), .B(\key_mem[9][55] ), .C(
        \key_mem[10][55] ), .D(\key_mem[11][55] ), .S0(n1381), .S1(n1311), .Y(
        n391) );
  MXI4X1 U5236 ( .A(\key_mem[8][21] ), .B(\key_mem[9][21] ), .C(
        \key_mem[10][21] ), .D(\key_mem[11][21] ), .S0(n1409), .S1(n1294), .Y(
        n207) );
  MXI4X1 U5237 ( .A(\key_mem[8][116] ), .B(\key_mem[9][116] ), .C(
        \key_mem[10][116] ), .D(\key_mem[11][116] ), .S0(n1391), .S1(n1301), 
        .Y(n1159) );
  MXI4X1 U5238 ( .A(\key_mem[8][84] ), .B(\key_mem[9][84] ), .C(
        \key_mem[10][84] ), .D(\key_mem[11][84] ), .S0(n1401), .S1(n1322), .Y(
        n536) );
  MXI4X1 U5239 ( .A(\key_mem[8][20] ), .B(\key_mem[9][20] ), .C(
        \key_mem[10][20] ), .D(\key_mem[11][20] ), .S0(n1408), .S1(n1293), .Y(
        n202) );
  MXI4X1 U5240 ( .A(\key_mem[8][115] ), .B(\key_mem[9][115] ), .C(
        \key_mem[10][115] ), .D(\key_mem[11][115] ), .S0(n1392), .S1(n1310), 
        .Y(n1139) );
  MXI4X1 U5241 ( .A(\key_mem[8][83] ), .B(\key_mem[9][83] ), .C(
        \key_mem[10][83] ), .D(\key_mem[11][83] ), .S0(n1401), .S1(n1322), .Y(
        n531) );
  MXI4X1 U5242 ( .A(\key_mem[8][114] ), .B(\key_mem[9][114] ), .C(
        \key_mem[10][114] ), .D(\key_mem[11][114] ), .S0(n1392), .S1(n1311), 
        .Y(n1125) );
  MXI4X1 U5243 ( .A(\key_mem[8][82] ), .B(\key_mem[9][82] ), .C(
        \key_mem[10][82] ), .D(\key_mem[11][82] ), .S0(n1402), .S1(n1322), .Y(
        n526) );
  MXI4X1 U5244 ( .A(\key_mem[8][18] ), .B(\key_mem[9][18] ), .C(
        \key_mem[10][18] ), .D(\key_mem[11][18] ), .S0(n1408), .S1(n1306), .Y(
        n168) );
  MXI4X1 U5245 ( .A(\key_mem[8][81] ), .B(\key_mem[9][81] ), .C(
        \key_mem[10][81] ), .D(\key_mem[11][81] ), .S0(n1402), .S1(n1321), .Y(
        n521) );
  MXI4X1 U5246 ( .A(\key_mem[8][17] ), .B(\key_mem[9][17] ), .C(
        \key_mem[10][17] ), .D(\key_mem[11][17] ), .S0(n1407), .S1(n1307), .Y(
        n163) );
  MXI4X1 U5247 ( .A(\key_mem[8][113] ), .B(\key_mem[9][113] ), .C(
        \key_mem[10][113] ), .D(\key_mem[11][113] ), .S0(n1392), .S1(n1313), 
        .Y(n1108) );
  MXI4X1 U5248 ( .A(\key_mem[8][80] ), .B(\key_mem[9][80] ), .C(
        \key_mem[10][80] ), .D(\key_mem[11][80] ), .S0(n1381), .S1(n1321), .Y(
        n516) );
  MXI4X1 U5249 ( .A(\key_mem[8][23] ), .B(\key_mem[9][23] ), .C(
        \key_mem[10][23] ), .D(\key_mem[11][23] ), .S0(n1409), .S1(n1295), .Y(
        n217) );
  MXI4X1 U5250 ( .A(\key_mem[8][118] ), .B(\key_mem[9][118] ), .C(
        \key_mem[10][118] ), .D(\key_mem[11][118] ), .S0(n1391), .S1(n1347), 
        .Y(n1180) );
  MXI4X1 U5251 ( .A(\key_mem[8][85] ), .B(\key_mem[9][85] ), .C(
        \key_mem[10][85] ), .D(\key_mem[11][85] ), .S0(n1401), .S1(n1323), .Y(
        n541) );
  MXI4X1 U5252 ( .A(\key_mem[8][53] ), .B(\key_mem[9][53] ), .C(
        \key_mem[10][53] ), .D(\key_mem[11][53] ), .S0(n1411), .S1(n1311), .Y(
        n381) );
  MXI4X1 U5253 ( .A(\key_mem[8][16] ), .B(\key_mem[9][16] ), .C(
        \key_mem[10][16] ), .D(\key_mem[11][16] ), .S0(n1407), .S1(n1330), .Y(
        n158) );
  MXI4X1 U5254 ( .A(\key_mem[8][117] ), .B(\key_mem[9][117] ), .C(
        \key_mem[10][117] ), .D(\key_mem[11][117] ), .S0(n1391), .S1(n1299), 
        .Y(n1171) );
  MXI4X1 U5255 ( .A(\key_mem[8][45] ), .B(\key_mem[9][45] ), .C(
        \key_mem[10][45] ), .D(\key_mem[11][45] ), .S0(n1413), .S1(n1305), .Y(
        n341) );
  MXI4X1 U5256 ( .A(\key_mem[8][109] ), .B(\key_mem[9][109] ), .C(
        \key_mem[10][109] ), .D(\key_mem[11][109] ), .S0(n1394), .S1(n1319), 
        .Y(n1027) );
  MXI4X1 U5257 ( .A(\key_mem[8][86] ), .B(\key_mem[9][86] ), .C(
        \key_mem[10][86] ), .D(\key_mem[11][86] ), .S0(n1401), .S1(n1323), .Y(
        n546) );
  MXI4X1 U5258 ( .A(\key_mem[8][54] ), .B(\key_mem[9][54] ), .C(
        \key_mem[10][54] ), .D(\key_mem[11][54] ), .S0(n1411), .S1(n1311), .Y(
        n386) );
  MXI4X1 U5259 ( .A(\key_mem[8][110] ), .B(\key_mem[9][110] ), .C(
        \key_mem[10][110] ), .D(\key_mem[11][110] ), .S0(n1393), .S1(n1317), 
        .Y(n1048) );
  MXI4X1 U5260 ( .A(\key_mem[8][46] ), .B(\key_mem[9][46] ), .C(
        \key_mem[10][46] ), .D(\key_mem[11][46] ), .S0(n1413), .S1(n1306), .Y(
        n346) );
  MXI4X1 U5261 ( .A(\key_mem[8][22] ), .B(\key_mem[9][22] ), .C(
        \key_mem[10][22] ), .D(\key_mem[11][22] ), .S0(n1409), .S1(n1303), .Y(
        n212) );
  MXI4X1 U5262 ( .A(\key_mem[8][78] ), .B(\key_mem[9][78] ), .C(
        \key_mem[10][78] ), .D(\key_mem[11][78] ), .S0(n1383), .S1(n1320), .Y(
        n506) );
  MXI4X1 U5263 ( .A(\key_mem[8][14] ), .B(\key_mem[9][14] ), .C(
        \key_mem[10][14] ), .D(\key_mem[11][14] ), .S0(n1406), .S1(n1329), .Y(
        n148) );
  MXI4X1 U5264 ( .A(\key_mem[8][77] ), .B(\key_mem[9][77] ), .C(
        \key_mem[10][77] ), .D(\key_mem[11][77] ), .S0(n1382), .S1(n1320), .Y(
        n501) );
  MXI4X1 U5265 ( .A(\key_mem[8][13] ), .B(\key_mem[9][13] ), .C(
        \key_mem[10][13] ), .D(\key_mem[11][13] ), .S0(n1406), .S1(n1329), .Y(
        n143) );
  MXI4X1 U5266 ( .A(\key_mem[8][12] ), .B(\key_mem[9][12] ), .C(
        \key_mem[10][12] ), .D(\key_mem[11][12] ), .S0(n1406), .S1(n1329), .Y(
        n138) );
  MXI4X1 U5267 ( .A(\key_mem[8][10] ), .B(\key_mem[9][10] ), .C(
        \key_mem[10][10] ), .D(\key_mem[11][10] ), .S0(n1405), .S1(n1328), .Y(
        n128) );
  MXI4X1 U5268 ( .A(\key_mem[8][9] ), .B(\key_mem[9][9] ), .C(\key_mem[10][9] ), .D(\key_mem[11][9] ), .S0(n1405), .S1(n1328), .Y(n123) );
  MXI4X1 U5269 ( .A(\key_mem[8][72] ), .B(\key_mem[9][72] ), .C(
        \key_mem[10][72] ), .D(\key_mem[11][72] ), .S0(n1385), .S1(n1318), .Y(
        n476) );
  MXI4X1 U5270 ( .A(\key_mem[8][8] ), .B(\key_mem[9][8] ), .C(\key_mem[10][8] ), .D(\key_mem[11][8] ), .S0(n1405), .S1(n1294), .Y(n118) );
  MXI4X1 U5271 ( .A(\key_mem[8][112] ), .B(\key_mem[9][112] ), .C(
        \key_mem[10][112] ), .D(\key_mem[11][112] ), .S0(n1393), .S1(n1314), 
        .Y(n1088) );
  MXI4X1 U5272 ( .A(\key_mem[8][47] ), .B(\key_mem[9][47] ), .C(
        \key_mem[10][47] ), .D(\key_mem[11][47] ), .S0(n1413), .S1(n1307), .Y(
        n351) );
  MXI4X1 U5273 ( .A(\key_mem[8][71] ), .B(\key_mem[9][71] ), .C(
        \key_mem[10][71] ), .D(\key_mem[11][71] ), .S0(n1386), .S1(n1317), .Y(
        n471) );
  MXI4X1 U5274 ( .A(\key_mem[8][15] ), .B(\key_mem[9][15] ), .C(
        \key_mem[10][15] ), .D(\key_mem[11][15] ), .S0(n1407), .S1(n1330), .Y(
        n153) );
  MXI4X1 U5275 ( .A(\key_mem[8][39] ), .B(\key_mem[9][39] ), .C(
        \key_mem[10][39] ), .D(\key_mem[11][39] ), .S0(n1415), .S1(n1297), .Y(
        n311) );
  MXI4X1 U5276 ( .A(\key_mem[8][111] ), .B(\key_mem[9][111] ), .C(
        \key_mem[10][111] ), .D(\key_mem[11][111] ), .S0(n1393), .S1(n1316), 
        .Y(n1068) );
  MXI4X1 U5277 ( .A(\key_mem[8][7] ), .B(\key_mem[9][7] ), .C(\key_mem[10][7] ), .D(\key_mem[11][7] ), .S0(n1404), .S1(n1303), .Y(n113) );
  MXI4X1 U5278 ( .A(\key_mem[8][79] ), .B(\key_mem[9][79] ), .C(
        \key_mem[10][79] ), .D(\key_mem[11][79] ), .S0(n1381), .S1(n1321), .Y(
        n511) );
  MXI4X1 U5279 ( .A(\key_mem[8][103] ), .B(\key_mem[9][103] ), .C(
        \key_mem[10][103] ), .D(\key_mem[11][103] ), .S0(n1395), .S1(n1303), 
        .Y(n956) );
  MXI4X1 U5280 ( .A(\key_mem[8][6] ), .B(\key_mem[9][6] ), .C(\key_mem[10][6] ), .D(\key_mem[11][6] ), .S0(n1404), .S1(n1304), .Y(n108) );
  MXI4X1 U5281 ( .A(\key_mem[8][38] ), .B(\key_mem[9][38] ), .C(
        \key_mem[10][38] ), .D(\key_mem[11][38] ), .S0(n1415), .S1(n1297), .Y(
        n306) );
  MXI4X1 U5282 ( .A(\key_mem[8][70] ), .B(\key_mem[9][70] ), .C(
        \key_mem[10][70] ), .D(\key_mem[11][70] ), .S0(n1383), .S1(n1317), .Y(
        n466) );
  MXI4X1 U5283 ( .A(\key_mem[8][102] ), .B(\key_mem[9][102] ), .C(
        \key_mem[10][102] ), .D(\key_mem[11][102] ), .S0(n1396), .S1(n1333), 
        .Y(n947) );
  MXI4X1 U5284 ( .A(\key_mem[8][5] ), .B(\key_mem[9][5] ), .C(\key_mem[10][5] ), .D(\key_mem[11][5] ), .S0(n1404), .S1(n1305), .Y(n103) );
  MXI4X1 U5285 ( .A(\key_mem[8][37] ), .B(\key_mem[9][37] ), .C(
        \key_mem[10][37] ), .D(\key_mem[11][37] ), .S0(n1353), .S1(n1297), .Y(
        n301) );
  MXI4X1 U5286 ( .A(\key_mem[8][69] ), .B(\key_mem[9][69] ), .C(
        \key_mem[10][69] ), .D(\key_mem[11][69] ), .S0(n1387), .S1(n1317), .Y(
        n461) );
  MXI4X1 U5287 ( .A(\key_mem[8][101] ), .B(\key_mem[9][101] ), .C(
        \key_mem[10][101] ), .D(\key_mem[11][101] ), .S0(n1396), .S1(n1327), 
        .Y(n936) );
  MXI4X1 U5288 ( .A(\key_mem[8][4] ), .B(\key_mem[9][4] ), .C(\key_mem[10][4] ), .D(\key_mem[11][4] ), .S0(n1403), .S1(n1307), .Y(n98) );
  MXI4X1 U5289 ( .A(\key_mem[8][36] ), .B(\key_mem[9][36] ), .C(
        \key_mem[10][36] ), .D(\key_mem[11][36] ), .S0(N31), .S1(n1309), .Y(
        n292) );
  MXI4X1 U5290 ( .A(\key_mem[8][68] ), .B(\key_mem[9][68] ), .C(
        \key_mem[10][68] ), .D(\key_mem[11][68] ), .S0(n1387), .S1(n1316), .Y(
        n456) );
  MXI4X1 U5291 ( .A(\key_mem[8][44] ), .B(\key_mem[9][44] ), .C(
        \key_mem[10][44] ), .D(\key_mem[11][44] ), .S0(n1414), .S1(n1296), .Y(
        n336) );
  MXI4X1 U5292 ( .A(\key_mem[8][108] ), .B(\key_mem[9][108] ), .C(
        \key_mem[10][108] ), .D(\key_mem[11][108] ), .S0(n1394), .S1(n1320), 
        .Y(n1007) );
  MXI4X1 U5293 ( .A(\key_mem[8][3] ), .B(\key_mem[9][3] ), .C(\key_mem[10][3] ), .D(\key_mem[11][3] ), .S0(n1403), .S1(n1307), .Y(n93) );
  MXI4X1 U5294 ( .A(\key_mem[8][67] ), .B(\key_mem[9][67] ), .C(
        \key_mem[10][67] ), .D(\key_mem[11][67] ), .S0(n1387), .S1(n1316), .Y(
        n451) );
  MXI4X1 U5295 ( .A(\key_mem[8][43] ), .B(\key_mem[9][43] ), .C(
        \key_mem[10][43] ), .D(\key_mem[11][43] ), .S0(n1414), .S1(n1303), .Y(
        n331) );
  MXI4X1 U5296 ( .A(\key_mem[8][42] ), .B(\key_mem[9][42] ), .C(
        \key_mem[10][42] ), .D(\key_mem[11][42] ), .S0(n1414), .S1(n1295), .Y(
        n326) );
  MXI4X1 U5297 ( .A(\key_mem[8][106] ), .B(\key_mem[9][106] ), .C(
        \key_mem[10][106] ), .D(\key_mem[11][106] ), .S0(n1394), .S1(n1323), 
        .Y(n987) );
  MXI4X1 U5298 ( .A(\key_mem[8][2] ), .B(\key_mem[9][2] ), .C(\key_mem[10][2] ), .D(\key_mem[11][2] ), .S0(n1403), .S1(n1300), .Y(n88) );
  MXI4X1 U5299 ( .A(\key_mem[8][34] ), .B(\key_mem[9][34] ), .C(
        \key_mem[10][34] ), .D(\key_mem[11][34] ), .S0(n1363), .S1(n1331), .Y(
        n272) );
  MXI4X1 U5300 ( .A(\key_mem[8][66] ), .B(\key_mem[9][66] ), .C(
        \key_mem[10][66] ), .D(\key_mem[11][66] ), .S0(n1388), .S1(n1316), .Y(
        n446) );
  MXI4X1 U5301 ( .A(\key_mem[8][1] ), .B(\key_mem[9][1] ), .C(\key_mem[10][1] ), .D(\key_mem[11][1] ), .S0(n1403), .S1(n1306), .Y(n83) );
  MXI4X1 U5302 ( .A(\key_mem[8][33] ), .B(\key_mem[9][33] ), .C(
        \key_mem[10][33] ), .D(\key_mem[11][33] ), .S0(n1353), .S1(n1332), .Y(
        n267) );
  MXI4X1 U5303 ( .A(\key_mem[8][65] ), .B(\key_mem[9][65] ), .C(
        \key_mem[10][65] ), .D(\key_mem[11][65] ), .S0(n1388), .S1(n1315), .Y(
        n441) );
  MXI4X1 U5304 ( .A(\key_mem[8][41] ), .B(\key_mem[9][41] ), .C(
        \key_mem[10][41] ), .D(\key_mem[11][41] ), .S0(n1414), .S1(n1297), .Y(
        n321) );
  MXI4X1 U5305 ( .A(\key_mem[8][105] ), .B(\key_mem[9][105] ), .C(
        \key_mem[10][105] ), .D(\key_mem[11][105] ), .S0(n1395), .S1(n1325), 
        .Y(n976) );
  MXI4X1 U5306 ( .A(\key_mem[8][40] ), .B(\key_mem[9][40] ), .C(
        \key_mem[10][40] ), .D(\key_mem[11][40] ), .S0(n1415), .S1(n1296), .Y(
        n316) );
  MXI4X1 U5307 ( .A(\key_mem[8][104] ), .B(\key_mem[9][104] ), .C(
        \key_mem[10][104] ), .D(\key_mem[11][104] ), .S0(n1395), .S1(n1326), 
        .Y(n967) );
  MXI4X1 U5308 ( .A(\key_mem[8][0] ), .B(\key_mem[9][0] ), .C(\key_mem[10][0] ), .D(\key_mem[11][0] ), .S0(n1402), .S1(n1327), .Y(n78) );
  MXI4X1 U5309 ( .A(\key_mem[8][32] ), .B(\key_mem[9][32] ), .C(
        \key_mem[10][32] ), .D(\key_mem[11][32] ), .S0(n1353), .S1(n1331), .Y(
        n262) );
  MXI4X1 U5310 ( .A(\key_mem[8][62] ), .B(\key_mem[9][62] ), .C(
        \key_mem[10][62] ), .D(\key_mem[11][62] ), .S0(n1385), .S1(n1314), .Y(
        n426) );
  MXI4X1 U5311 ( .A(\key_mem[8][29] ), .B(\key_mem[9][29] ), .C(
        \key_mem[10][29] ), .D(\key_mem[11][29] ), .S0(n1362), .S1(n1333), .Y(
        n247) );
  MXI4X1 U5312 ( .A(\key_mem[8][52] ), .B(\key_mem[9][52] ), .C(
        \key_mem[10][52] ), .D(\key_mem[11][52] ), .S0(n1411), .S1(n1310), .Y(
        n376) );
  MXI4X1 U5313 ( .A(\key_mem[8][28] ), .B(\key_mem[9][28] ), .C(
        \key_mem[10][28] ), .D(\key_mem[11][28] ), .S0(n1357), .S1(n1333), .Y(
        n242) );
  MXI4X1 U5314 ( .A(\key_mem[8][51] ), .B(\key_mem[9][51] ), .C(
        \key_mem[10][51] ), .D(\key_mem[11][51] ), .S0(n1411), .S1(n1310), .Y(
        n371) );
  MXI4X1 U5315 ( .A(\key_mem[8][27] ), .B(\key_mem[9][27] ), .C(
        \key_mem[10][27] ), .D(\key_mem[11][27] ), .S0(n1410), .S1(n1334), .Y(
        n237) );
  MXI4X1 U5316 ( .A(\key_mem[8][26] ), .B(\key_mem[9][26] ), .C(
        \key_mem[10][26] ), .D(\key_mem[11][26] ), .S0(n1410), .S1(n1309), .Y(
        n232) );
  MXI4X1 U5317 ( .A(\key_mem[8][25] ), .B(\key_mem[9][25] ), .C(
        \key_mem[10][25] ), .D(\key_mem[11][25] ), .S0(n1410), .S1(n1301), .Y(
        n227) );
  MXI4X1 U5318 ( .A(\key_mem[8][56] ), .B(\key_mem[9][56] ), .C(
        \key_mem[10][56] ), .D(\key_mem[11][56] ), .S0(n1381), .S1(n1312), .Y(
        n396) );
  MXI4X1 U5319 ( .A(\key_mem[8][61] ), .B(\key_mem[9][61] ), .C(
        \key_mem[10][61] ), .D(\key_mem[11][61] ), .S0(n1384), .S1(n1314), .Y(
        n421) );
  MXI4X1 U5320 ( .A(\key_mem[8][60] ), .B(\key_mem[9][60] ), .C(
        \key_mem[10][60] ), .D(\key_mem[11][60] ), .S0(n1384), .S1(n1313), .Y(
        n416) );
  MXI4X1 U5321 ( .A(\key_mem[8][59] ), .B(\key_mem[9][59] ), .C(
        \key_mem[10][59] ), .D(\key_mem[11][59] ), .S0(n1383), .S1(n1313), .Y(
        n411) );
  MXI4X1 U5322 ( .A(\key_mem[8][58] ), .B(\key_mem[9][58] ), .C(
        \key_mem[10][58] ), .D(\key_mem[11][58] ), .S0(n1382), .S1(n1313), .Y(
        n406) );
  MXI4X1 U5323 ( .A(\key_mem[8][57] ), .B(\key_mem[9][57] ), .C(
        \key_mem[10][57] ), .D(\key_mem[11][57] ), .S0(n1381), .S1(n1312), .Y(
        n401) );
  MXI4X1 U5324 ( .A(\key_mem[8][24] ), .B(\key_mem[9][24] ), .C(
        \key_mem[10][24] ), .D(\key_mem[11][24] ), .S0(n1409), .S1(n1294), .Y(
        n222) );
  MXI4X1 U5325 ( .A(\key_mem[8][31] ), .B(\key_mem[9][31] ), .C(
        \key_mem[10][31] ), .D(\key_mem[11][31] ), .S0(n1349), .S1(n1331), .Y(
        n257) );
  MXI4X1 U5326 ( .A(\key_mem[8][30] ), .B(\key_mem[9][30] ), .C(
        \key_mem[10][30] ), .D(\key_mem[11][30] ), .S0(n1364), .S1(n1333), .Y(
        n252) );
  MXI4X1 U5327 ( .A(\key_mem[8][126] ), .B(\key_mem[9][126] ), .C(
        \key_mem[10][126] ), .D(\key_mem[11][126] ), .S0(n1388), .S1(n1304), 
        .Y(n1257) );
  MXI4X1 U5328 ( .A(\key_mem[8][125] ), .B(\key_mem[9][125] ), .C(
        \key_mem[10][125] ), .D(\key_mem[11][125] ), .S0(n1389), .S1(n1328), 
        .Y(n1251) );
  MXI4X1 U5329 ( .A(\key_mem[8][124] ), .B(\key_mem[9][124] ), .C(
        \key_mem[10][124] ), .D(\key_mem[11][124] ), .S0(n1389), .S1(n1329), 
        .Y(n1240) );
  MXI4X1 U5330 ( .A(\key_mem[8][123] ), .B(\key_mem[9][123] ), .C(
        \key_mem[10][123] ), .D(\key_mem[11][123] ), .S0(n1389), .S1(n1302), 
        .Y(n1231) );
  MXI4X1 U5331 ( .A(\key_mem[8][122] ), .B(\key_mem[9][122] ), .C(
        \key_mem[10][122] ), .D(\key_mem[11][122] ), .S0(n1390), .S1(n1306), 
        .Y(n1220) );
  MXI4X1 U5332 ( .A(\key_mem[8][121] ), .B(\key_mem[9][121] ), .C(
        \key_mem[10][121] ), .D(\key_mem[11][121] ), .S0(n1390), .S1(n1303), 
        .Y(n1211) );
  MXI4X1 U5333 ( .A(\key_mem[8][120] ), .B(\key_mem[9][120] ), .C(
        \key_mem[10][120] ), .D(\key_mem[11][120] ), .S0(n1390), .S1(n1332), 
        .Y(n1200) );
  MXI4X1 U5334 ( .A(\key_mem[8][127] ), .B(\key_mem[9][127] ), .C(
        \key_mem[10][127] ), .D(\key_mem[11][127] ), .S0(n1388), .S1(n1298), 
        .Y(n1262) );
  MXI4X1 U5335 ( .A(\key_mem[8][94] ), .B(\key_mem[9][94] ), .C(
        \key_mem[10][94] ), .D(\key_mem[11][94] ), .S0(n1398), .S1(n1326), .Y(
        n586) );
  MXI4X1 U5336 ( .A(\key_mem[8][93] ), .B(\key_mem[9][93] ), .C(
        \key_mem[10][93] ), .D(\key_mem[11][93] ), .S0(n1398), .S1(n1326), .Y(
        n581) );
  MXI4X1 U5337 ( .A(\key_mem[8][92] ), .B(\key_mem[9][92] ), .C(
        \key_mem[10][92] ), .D(\key_mem[11][92] ), .S0(n1399), .S1(n1325), .Y(
        n576) );
  MXI4X1 U5338 ( .A(\key_mem[8][91] ), .B(\key_mem[9][91] ), .C(
        \key_mem[10][91] ), .D(\key_mem[11][91] ), .S0(n1399), .S1(n1325), .Y(
        n571) );
  MXI4X1 U5339 ( .A(\key_mem[8][90] ), .B(\key_mem[9][90] ), .C(
        \key_mem[10][90] ), .D(\key_mem[11][90] ), .S0(n1399), .S1(n1325), .Y(
        n566) );
  MXI4X1 U5340 ( .A(\key_mem[8][89] ), .B(\key_mem[9][89] ), .C(
        \key_mem[10][89] ), .D(\key_mem[11][89] ), .S0(n1400), .S1(n1324), .Y(
        n561) );
  MXI4X1 U5341 ( .A(\key_mem[8][88] ), .B(\key_mem[9][88] ), .C(
        \key_mem[10][88] ), .D(\key_mem[11][88] ), .S0(n1400), .S1(n1324), .Y(
        n556) );
  MXI4X1 U5342 ( .A(\key_mem[8][95] ), .B(\key_mem[9][95] ), .C(
        \key_mem[10][95] ), .D(\key_mem[11][95] ), .S0(n1398), .S1(n1347), .Y(
        n721) );
  MXI4X1 U5343 ( .A(\key_mem[8][63] ), .B(\key_mem[9][63] ), .C(
        \key_mem[10][63] ), .D(\key_mem[11][63] ), .S0(n1386), .S1(n1314), .Y(
        n431) );
  MXI4X1 U5344 ( .A(\key_mem[8][76] ), .B(\key_mem[9][76] ), .C(
        \key_mem[10][76] ), .D(\key_mem[11][76] ), .S0(n1382), .S1(n1319), .Y(
        n496) );
  MXI4X1 U5345 ( .A(\key_mem[8][74] ), .B(\key_mem[9][74] ), .C(
        \key_mem[10][74] ), .D(\key_mem[11][74] ), .S0(n1384), .S1(n1319), .Y(
        n486) );
  MXI4X1 U5346 ( .A(\key_mem[8][73] ), .B(\key_mem[9][73] ), .C(
        \key_mem[10][73] ), .D(\key_mem[11][73] ), .S0(n1385), .S1(n1318), .Y(
        n481) );
  MXI4X1 U5347 ( .A(\key_mem[8][100] ), .B(\key_mem[9][100] ), .C(
        \key_mem[10][100] ), .D(\key_mem[11][100] ), .S0(n1396), .S1(N32), .Y(
        n927) );
  MXI4X1 U5348 ( .A(\key_mem[8][99] ), .B(\key_mem[9][99] ), .C(
        \key_mem[10][99] ), .D(\key_mem[11][99] ), .S0(n1397), .S1(N32), .Y(
        n916) );
  MXI4X1 U5349 ( .A(\key_mem[8][98] ), .B(\key_mem[9][98] ), .C(
        \key_mem[10][98] ), .D(\key_mem[11][98] ), .S0(n1397), .S1(n1348), .Y(
        n907) );
  MXI4X1 U5350 ( .A(\key_mem[8][97] ), .B(\key_mem[9][97] ), .C(
        \key_mem[10][97] ), .D(\key_mem[11][97] ), .S0(n1397), .S1(N32), .Y(
        n767) );
  MXI4X1 U5351 ( .A(\key_mem[8][64] ), .B(\key_mem[9][64] ), .C(
        \key_mem[10][64] ), .D(\key_mem[11][64] ), .S0(n1387), .S1(n1315), .Y(
        n436) );
  MXI4X1 U5352 ( .A(\key_mem[8][96] ), .B(\key_mem[9][96] ), .C(
        \key_mem[10][96] ), .D(\key_mem[11][96] ), .S0(n1398), .S1(n1348), .Y(
        n748) );
  MXI4X1 U5353 ( .A(\key_mem[8][50] ), .B(\key_mem[9][50] ), .C(
        \key_mem[10][50] ), .D(\key_mem[11][50] ), .S0(n1412), .S1(n1310), .Y(
        n366) );
  MXI4X1 U5354 ( .A(\key_mem[8][49] ), .B(\key_mem[9][49] ), .C(
        \key_mem[10][49] ), .D(\key_mem[11][49] ), .S0(n1412), .S1(n1299), .Y(
        n361) );
  NOR2BX1 U5355 ( .AN(\key_mem[14][48] ), .B(n1360), .Y(n354) );
  NAND3BXL U5356 ( .AN(n1424), .B(keylen), .C(n4594), .Y(n4591) );
  NAND3BX1 U5357 ( .AN(n4588), .B(round_ctr_reg[0]), .C(n5760), .Y(n5762) );
  NOR3X1 U5358 ( .A(round_ctr_reg[2]), .B(round_ctr_reg[3]), .C(
        round_ctr_reg[1]), .Y(n1721) );
  NAND2BX1 U5359 ( .AN(n3976), .B(n4596), .Y(n4600) );
  AO21XL U5360 ( .A0(n4595), .A1(keylen), .B0(n1424), .Y(n4596) );
  INVX1 U5361 ( .A(n4594), .Y(n4595) );
  MXI4X1 U5362 ( .A(n196), .B(n197), .C(n198), .D(n199), .S0(n1270), .S1(n1285), .Y(round_key[19]) );
  MXI3X1 U5363 ( .A(\key_mem[12][19] ), .B(\key_mem[13][19] ), .C(n195), .S0(
        n1369), .S1(n1338), .Y(n199) );
  MXI4X1 U5364 ( .A(\key_mem[4][19] ), .B(\key_mem[5][19] ), .C(
        \key_mem[6][19] ), .D(\key_mem[7][19] ), .S0(n1408), .S1(n1293), .Y(
        n198) );
  MXI4X1 U5365 ( .A(\key_mem[0][19] ), .B(\key_mem[1][19] ), .C(
        \key_mem[2][19] ), .D(\key_mem[3][19] ), .S0(n1408), .S1(n1295), .Y(
        n196) );
  MXI4X1 U5366 ( .A(n132), .B(n133), .C(n134), .D(n135), .S0(N34), .S1(n1284), 
        .Y(round_key[11]) );
  MXI3X1 U5367 ( .A(\key_mem[12][11] ), .B(\key_mem[13][11] ), .C(n131), .S0(
        n1370), .S1(n1337), .Y(n135) );
  MXI4X1 U5368 ( .A(\key_mem[4][11] ), .B(\key_mem[5][11] ), .C(
        \key_mem[6][11] ), .D(\key_mem[7][11] ), .S0(n1406), .S1(n1328), .Y(
        n134) );
  MXI4X1 U5369 ( .A(\key_mem[0][11] ), .B(\key_mem[1][11] ), .C(
        \key_mem[2][11] ), .D(\key_mem[3][11] ), .S0(n1406), .S1(n1328), .Y(
        n132) );
  MXI4X1 U5370 ( .A(n280), .B(n282), .C(n284), .D(n286), .S0(n1271), .S1(n1286), .Y(round_key[35]) );
  MXI4X1 U5371 ( .A(\key_mem[4][35] ), .B(\key_mem[5][35] ), .C(
        \key_mem[6][35] ), .D(\key_mem[7][35] ), .S0(n1356), .S1(n1298), .Y(
        n284) );
  MXI3X1 U5372 ( .A(\key_mem[12][35] ), .B(\key_mem[13][35] ), .C(n275), .S0(
        n1374), .S1(n1340), .Y(n286) );
  MXI4X1 U5373 ( .A(\key_mem[0][35] ), .B(\key_mem[1][35] ), .C(
        \key_mem[2][35] ), .D(\key_mem[3][35] ), .S0(n1351), .S1(n1301), .Y(
        n280) );
  MXI4X1 U5374 ( .A(n995), .B(n996), .C(n999), .D(n1000), .S0(n1274), .S1(
        n1282), .Y(round_key[107]) );
  MXI4X1 U5375 ( .A(\key_mem[4][107] ), .B(\key_mem[5][107] ), .C(
        \key_mem[6][107] ), .D(\key_mem[7][107] ), .S0(n1394), .S1(n1321), .Y(
        n999) );
  MXI3X1 U5376 ( .A(\key_mem[12][107] ), .B(\key_mem[13][107] ), .C(n992), 
        .S0(n1375), .S1(n1334), .Y(n1000) );
  MXI4X1 U5377 ( .A(\key_mem[0][107] ), .B(\key_mem[1][107] ), .C(
        \key_mem[2][107] ), .D(\key_mem[3][107] ), .S0(n1394), .S1(n1321), .Y(
        n995) );
  MXI4X1 U5378 ( .A(n490), .B(n491), .C(n492), .D(n493), .S0(n1267), .S1(n1280), .Y(round_key[75]) );
  MXI4X1 U5379 ( .A(\key_mem[4][75] ), .B(\key_mem[5][75] ), .C(
        \key_mem[6][75] ), .D(\key_mem[7][75] ), .S0(n1383), .S1(n1319), .Y(
        n492) );
  MXI3X1 U5380 ( .A(\key_mem[12][75] ), .B(\key_mem[13][75] ), .C(n489), .S0(
        n1371), .S1(n1344), .Y(n493) );
  MXI4X1 U5381 ( .A(\key_mem[0][75] ), .B(\key_mem[1][75] ), .C(
        \key_mem[2][75] ), .D(\key_mem[3][75] ), .S0(n1383), .S1(n1319), .Y(
        n490) );
  NAND2BX1 U5382 ( .AN(key_mem_ctrl_reg[0]), .B(key_mem_ctrl_reg[1]), .Y(n5763) );
  NOR2BX1 U5383 ( .AN(\key_mem[14][83] ), .B(n1349), .Y(n529) );
  NOR2BX1 U5384 ( .AN(\key_mem[14][19] ), .B(n1356), .Y(n195) );
  NOR2BX1 U5385 ( .AN(\key_mem[14][11] ), .B(n1365), .Y(n131) );
  NOR2BX1 U5386 ( .AN(\key_mem[14][3] ), .B(n1355), .Y(n91) );
  NOR2BX1 U5387 ( .AN(\key_mem[14][35] ), .B(n1416), .Y(n275) );
  NOR2BX1 U5388 ( .AN(\key_mem[14][67] ), .B(n1360), .Y(n449) );
  NOR2BX1 U5389 ( .AN(\key_mem[14][43] ), .B(n1362), .Y(n329) );
  NOR2BX1 U5390 ( .AN(\key_mem[14][107] ), .B(n1349), .Y(n992) );
  NOR2BX1 U5391 ( .AN(\key_mem[14][51] ), .B(n1349), .Y(n369) );
  NOR2BX1 U5392 ( .AN(\key_mem[14][123] ), .B(n1358), .Y(n1227) );
  NOR2BX1 U5393 ( .AN(\key_mem[14][75] ), .B(N31), .Y(n489) );
  NOR2BX1 U5394 ( .AN(\key_mem[14][99] ), .B(n1353), .Y(n912) );
  MXI4X1 U5395 ( .A(\key_mem[8][19] ), .B(\key_mem[9][19] ), .C(
        \key_mem[10][19] ), .D(\key_mem[11][19] ), .S0(n1408), .S1(n1300), .Y(
        n197) );
  MXI4X1 U5396 ( .A(\key_mem[8][11] ), .B(\key_mem[9][11] ), .C(
        \key_mem[10][11] ), .D(\key_mem[11][11] ), .S0(n1406), .S1(n1328), .Y(
        n133) );
  MXI4X1 U5397 ( .A(\key_mem[8][35] ), .B(\key_mem[9][35] ), .C(
        \key_mem[10][35] ), .D(\key_mem[11][35] ), .S0(n1352), .S1(n1309), .Y(
        n282) );
  MXI4X1 U5398 ( .A(\key_mem[8][107] ), .B(\key_mem[9][107] ), .C(
        \key_mem[10][107] ), .D(\key_mem[11][107] ), .S0(n1394), .S1(n1322), 
        .Y(n996) );
  MXI4X1 U5399 ( .A(\key_mem[8][75] ), .B(\key_mem[9][75] ), .C(
        \key_mem[10][75] ), .D(\key_mem[11][75] ), .S0(n1383), .S1(n1319), .Y(
        n491) );
  XOR2X1 U5400 ( .A(n5425), .B(prev_key0_reg[89]), .Y(n5446) );
  XOR2X1 U5401 ( .A(n5533), .B(prev_key0_reg[92]), .Y(n5554) );
  XOR2X1 U5402 ( .A(n5569), .B(prev_key0_reg[93]), .Y(n5590) );
  XOR2X1 U5403 ( .A(n5605), .B(prev_key0_reg[94]), .Y(n5626) );
  XOR2X1 U5404 ( .A(n5497), .B(prev_key0_reg[91]), .Y(n5518) );
  XOR2X1 U5405 ( .A(n5461), .B(prev_key0_reg[90]), .Y(n5482) );
  XOR2X1 U5406 ( .A(n5389), .B(prev_key0_reg[88]), .Y(n5410) );
  XOR2X1 U5407 ( .A(n5446), .B(prev_key0_reg[57]), .Y(n5436) );
  XOR2X1 U5408 ( .A(n5554), .B(prev_key0_reg[60]), .Y(n5544) );
  XOR2X1 U5409 ( .A(n5590), .B(prev_key0_reg[61]), .Y(n5580) );
  XOR2X1 U5410 ( .A(n5626), .B(prev_key0_reg[62]), .Y(n5616) );
  XOR2X1 U5411 ( .A(n5518), .B(prev_key0_reg[59]), .Y(n5508) );
  XOR2X1 U5412 ( .A(n5482), .B(prev_key0_reg[58]), .Y(n5472) );
  XOR2X1 U5413 ( .A(n5410), .B(prev_key0_reg[56]), .Y(n5400) );
  XOR2X1 U5414 ( .A(n5641), .B(prev_key0_reg[95]), .Y(n5664) );
  XOR2X1 U5415 ( .A(n4640), .B(n193), .Y(n4659) );
  XOR2X1 U5416 ( .A(n4672), .B(n192), .Y(n4691) );
  XOR2X1 U5417 ( .A(n4704), .B(n191), .Y(n4723) );
  XOR2X1 U5418 ( .A(n4768), .B(n189), .Y(n4787) );
  XOR2X1 U5419 ( .A(n4799), .B(n188), .Y(n4818) );
  XOR2X1 U5420 ( .A(n4831), .B(n187), .Y(n4850) );
  XOR2X1 U5421 ( .A(n4897), .B(n185), .Y(n4916) );
  XOR2X1 U5422 ( .A(n4930), .B(n184), .Y(n4949) );
  XOR2X1 U5423 ( .A(n4963), .B(n183), .Y(n4982) );
  XOR2X1 U5424 ( .A(n5029), .B(n181), .Y(n5048) );
  XOR2X1 U5425 ( .A(n5094), .B(n179), .Y(n5113) );
  XOR2X1 U5426 ( .A(n5127), .B(n178), .Y(n5146) );
  XOR2X1 U5427 ( .A(n5160), .B(n177), .Y(n5179) );
  XOR2X1 U5428 ( .A(n5193), .B(n176), .Y(n5212) );
  XOR2X1 U5429 ( .A(n5226), .B(n175), .Y(n5245) );
  XOR2X1 U5430 ( .A(n5292), .B(n173), .Y(n5311) );
  XOR2X1 U5431 ( .A(n5325), .B(n172), .Y(n5343) );
  XOR2X1 U5432 ( .A(n5357), .B(n171), .Y(n5376) );
  XOR2X1 U5433 ( .A(n5259), .B(n174), .Y(n5278) );
  XOR2X1 U5434 ( .A(n5062), .B(n180), .Y(n5080) );
  XOR2X1 U5435 ( .A(n4609), .B(n194), .Y(n4627) );
  XOR2X1 U5436 ( .A(n4736), .B(n190), .Y(n4755) );
  XOR2X1 U5437 ( .A(n4864), .B(n186), .Y(n4883) );
  XOR2X1 U5438 ( .A(n4996), .B(n182), .Y(n5015) );
  XOR2X1 U5439 ( .A(n5426), .B(prev_key1_reg[89]), .Y(n5434) );
  XOR2X1 U5440 ( .A(n5534), .B(prev_key1_reg[92]), .Y(n5542) );
  XOR2X1 U5441 ( .A(n5570), .B(prev_key1_reg[93]), .Y(n5578) );
  XOR2X1 U5442 ( .A(n5606), .B(prev_key1_reg[94]), .Y(n5614) );
  XOR2X1 U5443 ( .A(n5498), .B(prev_key1_reg[91]), .Y(n5506) );
  XOR2X1 U5444 ( .A(n5462), .B(prev_key1_reg[90]), .Y(n5470) );
  XOR2X1 U5445 ( .A(n5390), .B(prev_key1_reg[88]), .Y(n5398) );
  XOR2X1 U5446 ( .A(n4659), .B(prev_key0_reg[33]), .Y(n4648) );
  XOR2X1 U5447 ( .A(n4691), .B(prev_key0_reg[34]), .Y(n4680) );
  XOR2X1 U5448 ( .A(n4723), .B(prev_key0_reg[35]), .Y(n4712) );
  XOR2X1 U5449 ( .A(n4787), .B(prev_key0_reg[37]), .Y(n4776) );
  XOR2X1 U5450 ( .A(n4818), .B(prev_key0_reg[38]), .Y(n4807) );
  XOR2X1 U5451 ( .A(n4850), .B(prev_key0_reg[39]), .Y(n4839) );
  XOR2X1 U5452 ( .A(n4949), .B(prev_key0_reg[42]), .Y(n4938) );
  XOR2X1 U5453 ( .A(n4982), .B(prev_key0_reg[43]), .Y(n4971) );
  XOR2X1 U5454 ( .A(n5048), .B(prev_key0_reg[45]), .Y(n5037) );
  XOR2X1 U5455 ( .A(n5080), .B(prev_key0_reg[46]), .Y(n5069) );
  XOR2X1 U5456 ( .A(n5113), .B(prev_key0_reg[47]), .Y(n5102) );
  XOR2X1 U5457 ( .A(n5212), .B(prev_key0_reg[50]), .Y(n5201) );
  XOR2X1 U5458 ( .A(n5245), .B(prev_key0_reg[51]), .Y(n5234) );
  XOR2X1 U5459 ( .A(n5311), .B(prev_key0_reg[53]), .Y(n5300) );
  XOR2X1 U5460 ( .A(n5376), .B(prev_key0_reg[55]), .Y(n5365) );
  XOR2X1 U5461 ( .A(n4627), .B(prev_key0_reg[32]), .Y(n4617) );
  XOR2X1 U5462 ( .A(n4755), .B(prev_key0_reg[36]), .Y(n4744) );
  XOR2X1 U5463 ( .A(n4883), .B(prev_key0_reg[40]), .Y(n4872) );
  XOR2X1 U5464 ( .A(n5179), .B(prev_key0_reg[49]), .Y(n5168) );
  XOR3X1 U5465 ( .A(prev_key0_reg[25]), .B(prev_key0_reg[57]), .C(n5446), .Y(
        n5449) );
  XOR3X1 U5466 ( .A(prev_key0_reg[28]), .B(prev_key0_reg[60]), .C(n5554), .Y(
        n5557) );
  XOR3X1 U5467 ( .A(prev_key0_reg[29]), .B(prev_key0_reg[61]), .C(n5590), .Y(
        n5593) );
  XOR3X1 U5468 ( .A(prev_key0_reg[30]), .B(prev_key0_reg[62]), .C(n5626), .Y(
        n5629) );
  XOR3X1 U5469 ( .A(prev_key0_reg[27]), .B(prev_key0_reg[59]), .C(n5518), .Y(
        n5521) );
  XOR3X1 U5470 ( .A(prev_key0_reg[26]), .B(prev_key0_reg[58]), .C(n5482), .Y(
        n5485) );
  XOR3X1 U5471 ( .A(prev_key0_reg[24]), .B(prev_key0_reg[56]), .C(n5410), .Y(
        n5413) );
  OAI22XL U5472 ( .A0(n287), .A1(n1722), .B0(n1723), .B1(n1724), .Y(n3916) );
  XNOR2X1 U5473 ( .A(rcon_reg[3]), .B(rcon_reg[7]), .Y(n1724) );
  OAI22XL U5474 ( .A0(n283), .A1(n1722), .B0(n1723), .B1(n285), .Y(n3914) );
  OAI22XL U5475 ( .A0(n285), .A1(n1722), .B0(n1723), .B1(n287), .Y(n3915) );
  OAI22XL U5476 ( .A0(n293), .A1(n1722), .B0(n1723), .B1(n1727), .Y(n3919) );
  XOR2X1 U5477 ( .A(n295), .B(rcon_reg[7]), .Y(n1727) );
  XOR3X1 U5478 ( .A(prev_key0_reg[31]), .B(prev_key0_reg[63]), .C(n5664), .Y(
        n5666) );
  XOR3X1 U5479 ( .A(prev_key0_reg[1]), .B(prev_key0_reg[33]), .C(n4659), .Y(
        n4660) );
  XOR3X1 U5480 ( .A(prev_key0_reg[2]), .B(prev_key0_reg[34]), .C(n4691), .Y(
        n4692) );
  XOR3X1 U5481 ( .A(prev_key0_reg[3]), .B(prev_key0_reg[35]), .C(n4723), .Y(
        n4724) );
  XOR3X1 U5482 ( .A(prev_key0_reg[5]), .B(prev_key0_reg[37]), .C(n4787), .Y(
        n4788) );
  XOR3X1 U5483 ( .A(prev_key0_reg[6]), .B(prev_key0_reg[38]), .C(n4818), .Y(
        n4819) );
  XOR3X1 U5484 ( .A(prev_key0_reg[7]), .B(prev_key0_reg[39]), .C(n4850), .Y(
        n4851) );
  XOR3X1 U5485 ( .A(prev_key0_reg[10]), .B(prev_key0_reg[42]), .C(n4949), .Y(
        n4950) );
  XOR3X1 U5486 ( .A(prev_key0_reg[11]), .B(prev_key0_reg[43]), .C(n4982), .Y(
        n4983) );
  XOR3X1 U5487 ( .A(prev_key0_reg[13]), .B(prev_key0_reg[45]), .C(n5048), .Y(
        n5049) );
  XOR3X1 U5488 ( .A(prev_key0_reg[14]), .B(prev_key0_reg[46]), .C(n5080), .Y(
        n5081) );
  XOR3X1 U5489 ( .A(prev_key0_reg[15]), .B(prev_key0_reg[47]), .C(n5113), .Y(
        n5114) );
  XOR3X1 U5490 ( .A(prev_key0_reg[16]), .B(prev_key0_reg[48]), .C(n5146), .Y(
        n5147) );
  XOR3X1 U5491 ( .A(prev_key0_reg[18]), .B(prev_key0_reg[50]), .C(n5212), .Y(
        n5213) );
  XOR3X1 U5492 ( .A(prev_key0_reg[19]), .B(prev_key0_reg[51]), .C(n5245), .Y(
        n5246) );
  XOR3X1 U5493 ( .A(prev_key0_reg[21]), .B(prev_key0_reg[53]), .C(n5311), .Y(
        n5312) );
  XOR3X1 U5494 ( .A(prev_key0_reg[23]), .B(prev_key0_reg[55]), .C(n5376), .Y(
        n5377) );
  XOR3X1 U5495 ( .A(prev_key0_reg[17]), .B(prev_key0_reg[49]), .C(n5179), .Y(
        n5180) );
  XOR3X1 U5496 ( .A(prev_key0_reg[0]), .B(prev_key0_reg[32]), .C(n4627), .Y(
        n4628) );
  XOR3X1 U5497 ( .A(prev_key0_reg[4]), .B(prev_key0_reg[36]), .C(n4755), .Y(
        n4756) );
  XOR3X1 U5498 ( .A(prev_key0_reg[8]), .B(prev_key0_reg[40]), .C(n4883), .Y(
        n4884) );
  XOR3X1 U5499 ( .A(prev_key0_reg[9]), .B(prev_key0_reg[41]), .C(n4916), .Y(
        n4917) );
  XOR3X1 U5500 ( .A(prev_key0_reg[12]), .B(prev_key0_reg[44]), .C(n5015), .Y(
        n5016) );
  XOR3X1 U5501 ( .A(prev_key0_reg[20]), .B(prev_key0_reg[52]), .C(n5278), .Y(
        n5279) );
  XOR3X1 U5502 ( .A(prev_key0_reg[22]), .B(prev_key0_reg[54]), .C(n5343), .Y(
        n5344) );
  NOR2BX1 U5503 ( .AN(n1718), .B(n726), .Y(n1723) );
  OA21XL U5504 ( .A0(keylen), .A1(n1424), .B0(n3985), .Y(n1718) );
  OAI221XL U5505 ( .A0(n1723), .A1(n1725), .B0(n289), .B1(n1722), .C0(n1726), 
        .Y(n3917) );
  XNOR2X1 U5506 ( .A(rcon_reg[2]), .B(rcon_reg[7]), .Y(n1725) );
  OAI221XL U5507 ( .A0(n1723), .A1(n293), .B0(n291), .B1(n1722), .C0(n1726), 
        .Y(n3918) );
  OAI221XL U5508 ( .A0(n1723), .A1(n281), .B0(n295), .B1(n1722), .C0(n1726), 
        .Y(n3920) );
  OAI221XL U5509 ( .A0(n1723), .A1(n283), .B0(n281), .B1(n1722), .C0(n1726), 
        .Y(n3921) );
  INVX1 U5510 ( .A(prev_key0_reg[102]), .Y(n4799) );
  INVX1 U5511 ( .A(prev_key0_reg[96]), .Y(n4609) );
  INVX1 U5512 ( .A(prev_key0_reg[98]), .Y(n4672) );
  INVX1 U5513 ( .A(prev_key0_reg[99]), .Y(n4704) );
  INVX1 U5514 ( .A(prev_key0_reg[100]), .Y(n4736) );
  INVX1 U5515 ( .A(prev_key0_reg[101]), .Y(n4768) );
  INVX1 U5516 ( .A(prev_key0_reg[103]), .Y(n4831) );
  INVX1 U5517 ( .A(prev_key0_reg[104]), .Y(n4864) );
  INVX1 U5518 ( .A(prev_key0_reg[106]), .Y(n4930) );
  INVX1 U5519 ( .A(prev_key0_reg[107]), .Y(n4963) );
  INVX1 U5520 ( .A(prev_key0_reg[109]), .Y(n5029) );
  INVX1 U5521 ( .A(prev_key0_reg[111]), .Y(n5094) );
  INVX1 U5522 ( .A(prev_key0_reg[113]), .Y(n5160) );
  INVX1 U5523 ( .A(prev_key0_reg[114]), .Y(n5193) );
  INVX1 U5524 ( .A(prev_key0_reg[115]), .Y(n5226) );
  INVX1 U5525 ( .A(prev_key0_reg[117]), .Y(n5292) );
  INVX1 U5526 ( .A(prev_key0_reg[119]), .Y(n5357) );
  INVX1 U5527 ( .A(prev_key0_reg[121]), .Y(n5425) );
  INVX1 U5528 ( .A(prev_key0_reg[124]), .Y(n5533) );
  INVX1 U5529 ( .A(prev_key0_reg[125]), .Y(n5569) );
  INVX1 U5530 ( .A(prev_key0_reg[126]), .Y(n5605) );
  INVX1 U5531 ( .A(prev_key0_reg[123]), .Y(n5497) );
  INVX1 U5532 ( .A(prev_key0_reg[122]), .Y(n5461) );
  INVX1 U5533 ( .A(prev_key0_reg[120]), .Y(n5389) );
  INVX1 U5534 ( .A(prev_key0_reg[127]), .Y(n5641) );
  INVX1 U5535 ( .A(prev_key0_reg[97]), .Y(n4640) );
  INVX1 U5536 ( .A(prev_key0_reg[110]), .Y(n5062) );
  INVX1 U5537 ( .A(prev_key1_reg[121]), .Y(n5426) );
  INVX1 U5538 ( .A(prev_key1_reg[124]), .Y(n5534) );
  INVX1 U5539 ( .A(prev_key1_reg[125]), .Y(n5570) );
  INVX1 U5540 ( .A(prev_key1_reg[126]), .Y(n5606) );
  INVX1 U5541 ( .A(prev_key1_reg[123]), .Y(n5498) );
  INVX1 U5542 ( .A(prev_key1_reg[122]), .Y(n5462) );
  INVX1 U5543 ( .A(prev_key1_reg[120]), .Y(n5390) );
  NOR2X1 U5544 ( .A(n5763), .B(round_ctr_reg[0]), .Y(n723) );
  NOR2X1 U5545 ( .A(n279), .B(n1424), .Y(n726) );
  NOR2X1 U5546 ( .A(n277), .B(round_ctr_reg[1]), .Y(n728) );
  XOR2X1 U5547 ( .A(n5643), .B(prev_key1_reg[95]), .Y(n5651) );
  XOR2X1 U5548 ( .A(n5343), .B(prev_key0_reg[54]), .Y(n5333) );
  XOR2X1 U5549 ( .A(n5146), .B(prev_key0_reg[48]), .Y(n5135) );
  XOR2X1 U5550 ( .A(n5664), .B(prev_key0_reg[63]), .Y(n5652) );
  XOR2X1 U5551 ( .A(n4916), .B(prev_key0_reg[41]), .Y(n4905) );
  NAND4X1 U5552 ( .A(round_ctr_reg[3]), .B(round_ctr_reg[2]), .C(n723), .D(
        round_ctr_reg[1]), .Y(n740) );
  NOR3X1 U5553 ( .A(round_ctr_reg[2]), .B(round_ctr_reg[3]), .C(n278), .Y(n724) );
  XOR2X1 U5554 ( .A(n5278), .B(prev_key0_reg[52]), .Y(n5267) );
  NAND3X1 U5555 ( .A(n726), .B(round_ctr_reg[1]), .C(n734), .Y(n737) );
  NAND3X1 U5556 ( .A(n723), .B(round_ctr_reg[1]), .C(n734), .Y(n736) );
  OAI22XL U5557 ( .A0(n1731), .A1(n278), .B0(round_ctr_reg[1]), .B1(n1729), 
        .Y(n3924) );
  XOR2X1 U5558 ( .A(n5015), .B(prev_key0_reg[44]), .Y(n5004) );
  NAND3X1 U5559 ( .A(n723), .B(n278), .C(n734), .Y(n733) );
  NAND3X1 U5560 ( .A(n723), .B(n276), .C(n728), .Y(n727) );
  NAND3X1 U5561 ( .A(n728), .B(n726), .C(round_ctr_reg[3]), .Y(n739) );
  NAND3X1 U5562 ( .A(n728), .B(n723), .C(round_ctr_reg[3]), .Y(n738) );
  NAND3X1 U5563 ( .A(n726), .B(n278), .C(n734), .Y(n735) );
  NAND3X1 U5564 ( .A(n726), .B(n276), .C(n728), .Y(n729) );
  OR2X1 U5565 ( .A(n276), .B(round_ctr_reg[2]), .Y(n5764) );
  NAND3BX1 U5566 ( .AN(key_mem_ctrl_reg[1]), .B(n299), .C(init), .Y(n591) );
  NAND3X1 U5567 ( .A(round_ctr_reg[1]), .B(round_ctr_reg[2]), .C(n276), .Y(
        n731) );
  NAND4X1 U5568 ( .A(n75), .B(round_ctr_reg[3]), .C(round_ctr_reg[1]), .D(n279), .Y(n1734) );
  NAND2X1 U5569 ( .A(round_ctr_reg[0]), .B(n5760), .Y(n1729) );
  NAND2X1 U5570 ( .A(n298), .B(key_mem_ctrl_reg[0]), .Y(n1733) );
  OA21XL U5571 ( .A0(round_ctr_reg[0]), .A1(n5763), .B0(n1732), .Y(n1731) );
  OA21XL U5572 ( .A0(round_ctr_reg[1]), .A1(n1424), .B0(n1731), .Y(n1730) );
  OAI222XL U5573 ( .A0(n731), .A1(n1729), .B0(n5763), .B1(n5764), .C0(n1730), 
        .C1(n276), .Y(n3922) );
  OAI221XL U5574 ( .A0(n298), .A1(n1734), .B0(key_mem_ctrl_reg[1]), .B1(n5765), 
        .C0(n299), .Y(n1735) );
  INVX1 U5575 ( .A(init), .Y(n5765) );
  OAI32X1 U5576 ( .A0(n1729), .A1(round_ctr_reg[2]), .A2(n278), .B0(n1730), 
        .B1(n277), .Y(n3923) );
  OAI221XL U5577 ( .A0(n1424), .A1(n1734), .B0(n1735), .B1(n299), .C0(n591), 
        .Y(n3927) );
  OAI211X1 U5578 ( .A0(n1735), .A1(n298), .B0(n1733), .C0(n1424), .Y(n3926) );
  INVX1 U5579 ( .A(prev_key0_reg[118]), .Y(n5325) );
  INVX1 U5580 ( .A(prev_key0_reg[112]), .Y(n5127) );
  INVX1 U5581 ( .A(prev_key0_reg[116]), .Y(n5259) );
  INVX1 U5582 ( .A(prev_key0_reg[105]), .Y(n4897) );
  INVX1 U5583 ( .A(prev_key1_reg[127]), .Y(n5643) );
  INVX1 U5584 ( .A(prev_key0_reg[108]), .Y(n4996) );
  OAI21XL U5585 ( .A0(n298), .A1(n299), .B0(n590), .Y(n1737) );
  NAND2X1 U5586 ( .A(ready), .B(n591), .Y(n590) );
  INVX1 U5587 ( .A(key[54]), .Y(n5337) );
  INVX1 U5588 ( .A(key[78]), .Y(n5066) );
  INVX1 U5589 ( .A(key[200]), .Y(n5785) );
  INVX1 U5590 ( .A(key[176]), .Y(n5793) );
  INVX1 U5591 ( .A(key[137]), .Y(n5773) );
  INVX1 U5592 ( .A(key[140]), .Y(n5837) );
  INVX1 U5593 ( .A(key[144]), .Y(n5791) );
  INVX1 U5594 ( .A(key[145]), .Y(n5779) );
  INVX1 U5595 ( .A(key[169]), .Y(n5767) );
  INVX1 U5596 ( .A(key[172]), .Y(n5835) );
  INVX1 U5597 ( .A(key[177]), .Y(n5777) );
  INVX1 U5598 ( .A(key[180]), .Y(n5841) );
  INVX1 U5599 ( .A(key[201]), .Y(n5772) );
  INVX1 U5600 ( .A(key[204]), .Y(n5833) );
  INVX1 U5601 ( .A(key[208]), .Y(n5795) );
  INVX1 U5602 ( .A(key[214]), .Y(n5875) );
  INVX1 U5603 ( .A(key[206]), .Y(n5865) );
  INVX1 U5604 ( .A(key[132]), .Y(n5838) );
  INVX1 U5605 ( .A(key[136]), .Y(n5789) );
  INVX1 U5606 ( .A(key[168]), .Y(n5787) );
  INVX1 U5607 ( .A(key[192]), .Y(n5794) );
  INVX1 U5608 ( .A(key[196]), .Y(n5842) );
  INVX1 U5609 ( .A(key[236]), .Y(n5831) );
  INVX1 U5610 ( .A(key[153]), .Y(n5771) );
  INVX1 U5611 ( .A(key[185]), .Y(n5769) );
  INVX1 U5612 ( .A(key[217]), .Y(n5770) );
  INVX1 U5613 ( .A(key[249]), .Y(n5768) );
  INVX1 U5614 ( .A(key[156]), .Y(n5836) );
  INVX1 U5615 ( .A(key[188]), .Y(n5834) );
  INVX1 U5616 ( .A(key[220]), .Y(n5832) );
  INVX1 U5617 ( .A(key[252]), .Y(n5830) );
  INVX1 U5618 ( .A(key[157]), .Y(n5852) );
  INVX1 U5619 ( .A(key[189]), .Y(n5850) );
  INVX1 U5620 ( .A(key[221]), .Y(n5848) );
  INVX1 U5621 ( .A(key[253]), .Y(n5846) );
  INVX1 U5622 ( .A(key[158]), .Y(n5868) );
  INVX1 U5623 ( .A(key[190]), .Y(n5866) );
  INVX1 U5624 ( .A(key[222]), .Y(n5864) );
  INVX1 U5625 ( .A(key[254]), .Y(n5862) );
  INVX1 U5626 ( .A(key[155]), .Y(n5820) );
  INVX1 U5627 ( .A(key[187]), .Y(n5818) );
  INVX1 U5628 ( .A(key[219]), .Y(n5816) );
  INVX1 U5629 ( .A(key[251]), .Y(n5814) );
  INVX1 U5630 ( .A(key[154]), .Y(n5804) );
  INVX1 U5631 ( .A(key[186]), .Y(n5802) );
  INVX1 U5632 ( .A(key[218]), .Y(n5800) );
  INVX1 U5633 ( .A(key[250]), .Y(n5798) );
  INVX1 U5634 ( .A(key[152]), .Y(n5788) );
  INVX1 U5635 ( .A(key[184]), .Y(n5786) );
  INVX1 U5636 ( .A(key[216]), .Y(n5784) );
  INVX1 U5637 ( .A(key[248]), .Y(n5782) );
  INVX1 U5638 ( .A(key[159]), .Y(n5884) );
  INVX1 U5639 ( .A(key[191]), .Y(n5882) );
  INVX1 U5640 ( .A(key[223]), .Y(n5880) );
  INVX1 U5641 ( .A(key[255]), .Y(n5878) );
  INVX1 U5642 ( .A(key[128]), .Y(n5790) );
  INVX1 U5643 ( .A(key[129]), .Y(n5781) );
  INVX1 U5644 ( .A(key[130]), .Y(n5806) );
  INVX1 U5645 ( .A(key[131]), .Y(n5822) );
  INVX1 U5646 ( .A(key[133]), .Y(n5854) );
  INVX1 U5647 ( .A(key[134]), .Y(n5870) );
  INVX1 U5648 ( .A(key[135]), .Y(n5886) );
  INVX1 U5649 ( .A(key[138]), .Y(n5805) );
  INVX1 U5650 ( .A(key[139]), .Y(n5821) );
  INVX1 U5651 ( .A(key[141]), .Y(n5853) );
  INVX1 U5652 ( .A(key[142]), .Y(n5869) );
  INVX1 U5653 ( .A(key[143]), .Y(n5885) );
  INVX1 U5654 ( .A(key[146]), .Y(n5807) );
  INVX1 U5655 ( .A(key[147]), .Y(n5823) );
  INVX1 U5656 ( .A(key[148]), .Y(n5839) );
  INVX1 U5657 ( .A(key[149]), .Y(n5855) );
  INVX1 U5658 ( .A(key[150]), .Y(n5871) );
  INVX1 U5659 ( .A(key[151]), .Y(n5887) );
  INVX1 U5660 ( .A(key[160]), .Y(n5792) );
  INVX1 U5661 ( .A(key[161]), .Y(n5775) );
  INVX1 U5662 ( .A(key[162]), .Y(n5808) );
  INVX1 U5663 ( .A(key[163]), .Y(n5824) );
  INVX1 U5664 ( .A(key[164]), .Y(n5840) );
  INVX1 U5665 ( .A(key[165]), .Y(n5856) );
  INVX1 U5666 ( .A(key[166]), .Y(n5872) );
  INVX1 U5667 ( .A(key[167]), .Y(n5888) );
  INVX1 U5668 ( .A(key[170]), .Y(n5803) );
  INVX1 U5669 ( .A(key[171]), .Y(n5819) );
  INVX1 U5670 ( .A(key[173]), .Y(n5851) );
  INVX1 U5671 ( .A(key[174]), .Y(n5867) );
  INVX1 U5672 ( .A(key[175]), .Y(n5883) );
  INVX1 U5673 ( .A(key[178]), .Y(n5809) );
  INVX1 U5674 ( .A(key[179]), .Y(n5825) );
  INVX1 U5675 ( .A(key[181]), .Y(n5857) );
  INVX1 U5676 ( .A(key[182]), .Y(n5873) );
  INVX1 U5677 ( .A(key[183]), .Y(n5889) );
  INVX1 U5678 ( .A(key[193]), .Y(n5780) );
  INVX1 U5679 ( .A(key[194]), .Y(n5810) );
  INVX1 U5680 ( .A(key[195]), .Y(n5826) );
  INVX1 U5681 ( .A(key[197]), .Y(n5858) );
  INVX1 U5682 ( .A(key[198]), .Y(n5874) );
  INVX1 U5683 ( .A(key[199]), .Y(n5890) );
  INVX1 U5684 ( .A(key[202]), .Y(n5801) );
  INVX1 U5685 ( .A(key[203]), .Y(n5817) );
  INVX1 U5686 ( .A(key[205]), .Y(n5849) );
  INVX1 U5687 ( .A(key[207]), .Y(n5881) );
  INVX1 U5688 ( .A(key[209]), .Y(n5778) );
  INVX1 U5689 ( .A(key[210]), .Y(n5811) );
  INVX1 U5690 ( .A(key[211]), .Y(n5827) );
  INVX1 U5691 ( .A(key[212]), .Y(n5843) );
  INVX1 U5692 ( .A(key[213]), .Y(n5859) );
  INVX1 U5693 ( .A(key[215]), .Y(n5891) );
  INVX1 U5694 ( .A(key[224]), .Y(n5796) );
  INVX1 U5695 ( .A(key[225]), .Y(n5774) );
  INVX1 U5696 ( .A(key[226]), .Y(n5812) );
  INVX1 U5697 ( .A(key[227]), .Y(n5828) );
  INVX1 U5698 ( .A(key[228]), .Y(n5844) );
  INVX1 U5699 ( .A(key[229]), .Y(n5860) );
  INVX1 U5700 ( .A(key[230]), .Y(n5876) );
  INVX1 U5701 ( .A(key[231]), .Y(n5892) );
  INVX1 U5702 ( .A(key[232]), .Y(n5783) );
  INVX1 U5703 ( .A(key[233]), .Y(n5766) );
  INVX1 U5704 ( .A(key[234]), .Y(n5799) );
  INVX1 U5705 ( .A(key[235]), .Y(n5815) );
  INVX1 U5706 ( .A(key[237]), .Y(n5847) );
  INVX1 U5707 ( .A(key[238]), .Y(n5863) );
  INVX1 U5708 ( .A(key[239]), .Y(n5879) );
  INVX1 U5709 ( .A(key[240]), .Y(n5797) );
  INVX1 U5710 ( .A(key[241]), .Y(n5776) );
  INVX1 U5711 ( .A(key[242]), .Y(n5813) );
  INVX1 U5712 ( .A(key[243]), .Y(n5829) );
  INVX1 U5713 ( .A(key[244]), .Y(n5845) );
  INVX1 U5714 ( .A(key[245]), .Y(n5861) );
  INVX1 U5715 ( .A(key[246]), .Y(n5877) );
  INVX1 U5716 ( .A(key[247]), .Y(n5893) );
  MXI4X1 U5717 ( .A(\key_mem[0][48] ), .B(\key_mem[1][48] ), .C(
        \key_mem[2][48] ), .D(\key_mem[3][48] ), .S0(n1412), .S1(n1299), .Y(
        n355) );
  MXI4X1 U5718 ( .A(\key_mem[4][48] ), .B(\key_mem[5][48] ), .C(
        \key_mem[6][48] ), .D(\key_mem[7][48] ), .S0(n1412), .S1(n1293), .Y(
        n357) );
  MXI4X1 U5719 ( .A(\key_mem[8][48] ), .B(\key_mem[9][48] ), .C(
        \key_mem[10][48] ), .D(\key_mem[11][48] ), .S0(n1412), .S1(n1301), .Y(
        n356) );
  MXI3X1 U5720 ( .A(\key_mem[12][48] ), .B(\key_mem[13][48] ), .C(n354), .S0(
        n1379), .S1(n1341), .Y(n358) );
  INVX1 U5721 ( .A(n5728), .Y(n4909) );
  INVX1 U5722 ( .A(n5729), .Y(n4901) );
  INVXL U5723 ( .A(n4661), .Y(n1249) );
  INVXL U5724 ( .A(n4649), .Y(n1121) );
  INVXL U5725 ( .A(n4641), .Y(n993) );
  XOR2X1 U5726 ( .A(n4891), .B(prev_key0_reg[105]), .Y(n4895) );
  AO22XL U5727 ( .A0(sboxw[4]), .A1(n1618), .B0(n1604), .B1(n4757), .Y(n4758)
         );
  XNOR2X1 U5728 ( .A(prev_key0_reg[102]), .B(n5056), .Y(n1419) );
  XOR2X1 U5729 ( .A(n4628), .B(n4858), .Y(n1422) );
  INVXL U5730 ( .A(n5696), .Y(n5271) );
  AO22XL U5731 ( .A0(sboxw[12]), .A1(n1609), .B0(n1596), .B1(n5017), .Y(n5018)
         );
  INVXL U5732 ( .A(n5017), .Y(n1205) );
  AO22XL U5733 ( .A0(prev_key1_reg[44]), .A1(n1609), .B0(n1596), .B1(n5005), 
        .Y(n5006) );
  INVXL U5734 ( .A(n5005), .Y(n1077) );
  AO22XL U5735 ( .A0(prev_key1_reg[76]), .A1(n1618), .B0(n1605), .B1(n4997), 
        .Y(n4998) );
  INVXL U5736 ( .A(n4997), .Y(n949) );
  OAI2BB2XL U5737 ( .B0(n4603), .B1(n3), .A0N(prev_key1_reg[32]), .A1N(n1608), 
        .Y(n4618) );
  NAND2BX1 U5738 ( .AN(round_ctr_reg[0]), .B(n4592), .Y(n4593) );
  INVX1 U5739 ( .A(n5708), .Y(n5139) );
  INVX1 U5740 ( .A(n4865), .Y(n965) );
  INVXL U5741 ( .A(n837), .Y(n4859) );
  INVX1 U5742 ( .A(n5707), .Y(n5151) );
  INVX1 U5743 ( .A(n5719), .Y(n5008) );
  INVX1 U5744 ( .A(n5720), .Y(n5000) );
  INVXL U5745 ( .A(n4757), .Y(n1237) );
  INVXL U5746 ( .A(n4737), .Y(n981) );
  INVXL U5747 ( .A(n853), .Y(n4731) );
  INVXL U5748 ( .A(n5718), .Y(n5020) );
  INVXL U5749 ( .A(n5727), .Y(n4921) );
  AO22XL U5750 ( .A0(prev_key1_reg[78]), .A1(n1609), .B0(n1596), .B1(n5063), 
        .Y(n5064) );
  INVXL U5751 ( .A(n5063), .Y(n941) );
  AO22XL U5752 ( .A0(prev_key1_reg[64]), .A1(n1608), .B0(n1595), .B1(n4610), 
        .Y(n4611) );
  INVXL U5753 ( .A(n4610), .Y(n997) );
  AO22XL U5754 ( .A0(prev_key1_reg[110]), .A1(n1609), .B0(n1596), .B1(n5057), 
        .Y(n5058) );
  INVXL U5755 ( .A(n813), .Y(n5057) );
  AO22XL U5756 ( .A0(prev_key1_reg[108]), .A1(n1620), .B0(n1602), .B1(n4991), 
        .Y(n4992) );
  INVXL U5757 ( .A(n821), .Y(n4991) );
  INVXL U5758 ( .A(n5709), .Y(n5131) );
  AO22XL U5759 ( .A0(prev_key1_reg[97]), .A1(n1608), .B0(n1595), .B1(n4635), 
        .Y(n4636) );
  INVXL U5760 ( .A(n865), .Y(n4635) );
  AOI222XL U5761 ( .A0(n1707), .A1(n68), .B0(key[86]), .B1(n1682), .C0(n1702), 
        .C1(n5691), .Y(n910) );
  INVXL U5762 ( .A(n4745), .Y(n1109) );
  AO22XL U5763 ( .A0(sboxw[8]), .A1(n1617), .B0(n1605), .B1(n4885), .Y(n4886)
         );
  INVXL U5764 ( .A(n4885), .Y(n1221) );
  INVXL U5765 ( .A(n5690), .Y(n5348) );
  AOI222XL U5766 ( .A0(n1712), .A1(n74), .B0(key[22]), .B1(n1689), .C0(n1702), 
        .C1(n5690), .Y(n1166) );
  AOI222XL U5767 ( .A0(n1708), .A1(n11), .B0(key[72]), .B1(n1682), .C0(n1695), 
        .C1(n5732), .Y(n966) );
  INVXL U5768 ( .A(n5732), .Y(n4868) );
  AOI222XL U5769 ( .A0(n1711), .A1(n1095), .B0(key[40]), .B1(n1684), .C0(n1698), .C1(n5731), .Y(n1094) );
  AOI222XL U5770 ( .A0(n1714), .A1(n9), .B0(key[8]), .B1(n1685), .C0(n1699), 
        .C1(n5730), .Y(n1222) );
  AO22XL U5771 ( .A0(prev_key1_reg[40]), .A1(n1619), .B0(n1607), .B1(n4873), 
        .Y(n4874) );
  INVXL U5772 ( .A(n4873), .Y(n1093) );
  AO22XL U5773 ( .A0(prev_key1_reg[72]), .A1(n1619), .B0(n1603), .B1(n4865), 
        .Y(n4866) );
  AOI222XL U5774 ( .A0(n1711), .A1(n1071), .B0(key[46]), .B1(n1684), .C0(n1698), .C1(n5714), .Y(n1070) );
  INVXL U5775 ( .A(n5705), .Y(n5172) );
  AOI222XL U5776 ( .A0(n1713), .A1(n10), .B0(key[14]), .B1(n1687), .C0(n1699), 
        .C1(n5713), .Y(n1198) );
  AOI222XL U5777 ( .A0(n1707), .A1(n67), .B0(key[81]), .B1(n1682), .C0(n1703), 
        .C1(n5706), .Y(n930) );
  AOI222XL U5778 ( .A0(n1708), .A1(n31), .B0(key[73]), .B1(n1690), .C0(n1695), 
        .C1(n5729), .Y(n962) );
  AOI222XL U5779 ( .A0(n1707), .A1(n66), .B0(key[80]), .B1(n1682), .C0(n1699), 
        .C1(n5709), .Y(n934) );
  AOI222XL U5780 ( .A0(n1711), .A1(n1063), .B0(key[48]), .B1(n1683), .C0(n1698), .C1(n5708), .Y(n1062) );
  INVXL U5781 ( .A(n5697), .Y(n5263) );
  AOI222XL U5782 ( .A0(n1708), .A1(n69), .B0(key[76]), .B1(n1687), .C0(n1695), 
        .C1(n5720), .Y(n950) );
  AOI222XL U5783 ( .A0(n1710), .A1(n1047), .B0(key[52]), .B1(n1683), .C0(n1697), .C1(n5696), .Y(n1046) );
  AOI222XL U5784 ( .A0(n1711), .A1(n1091), .B0(key[41]), .B1(n1684), .C0(n1698), .C1(n5728), .Y(n1090) );
  AOI222XL U5785 ( .A0(n1711), .A1(n1079), .B0(key[44]), .B1(n1684), .C0(n1698), .C1(n5719), .Y(n1078) );
  AOI222XL U5786 ( .A0(n1710), .A1(n1059), .B0(key[49]), .B1(n1683), .C0(n1697), .C1(n5705), .Y(n1058) );
  INVXL U5787 ( .A(n5695), .Y(n5283) );
  AOI222XL U5788 ( .A0(n1713), .A1(n70), .B0(key[9]), .B1(n1689), .C0(n5758), 
        .C1(n5727), .Y(n1218) );
  AOI222XL U5789 ( .A0(n1713), .A1(n71), .B0(key[16]), .B1(n1687), .C0(n1702), 
        .C1(n5707), .Y(n1190) );
  AOI222XL U5790 ( .A0(n1714), .A1(n72), .B0(key[17]), .B1(n1685), .C0(n1703), 
        .C1(n5704), .Y(n1186) );
  AOI222XL U5791 ( .A0(n1712), .A1(n73), .B0(key[20]), .B1(n1686), .C0(n1702), 
        .C1(n5695), .Y(n1174) );
  INVX1 U5792 ( .A(n4575), .Y(n4370) );
  INVX1 U5793 ( .A(n4575), .Y(n4371) );
  INVX1 U5794 ( .A(n4575), .Y(n4372) );
  INVX1 U5795 ( .A(n4575), .Y(n4373) );
  INVX1 U5796 ( .A(n4575), .Y(n4374) );
  INVX1 U5797 ( .A(n4575), .Y(n4375) );
  INVX1 U5798 ( .A(n4575), .Y(n4376) );
  INVX1 U5799 ( .A(n4575), .Y(n4377) );
  INVX1 U5800 ( .A(n4575), .Y(n4378) );
  INVX1 U5801 ( .A(n4575), .Y(n4379) );
  INVX1 U5802 ( .A(n4574), .Y(n4380) );
  INVX1 U5803 ( .A(n4574), .Y(n4381) );
  INVX1 U5804 ( .A(n4574), .Y(n4382) );
  INVX1 U5805 ( .A(n4574), .Y(n4383) );
  INVX1 U5806 ( .A(n4574), .Y(n4384) );
  INVX1 U5807 ( .A(n4574), .Y(n4385) );
  INVX1 U5808 ( .A(n4574), .Y(n4386) );
  INVX1 U5809 ( .A(n4574), .Y(n4387) );
  INVX1 U5810 ( .A(n4574), .Y(n4388) );
  INVX1 U5811 ( .A(n4574), .Y(n4389) );
  INVX1 U5812 ( .A(n4573), .Y(n4390) );
  INVX1 U5813 ( .A(n4573), .Y(n4391) );
  INVX1 U5814 ( .A(n4573), .Y(n4392) );
  INVX1 U5815 ( .A(n4573), .Y(n4393) );
  INVX1 U5816 ( .A(n4573), .Y(n4394) );
  INVX1 U5817 ( .A(n4573), .Y(n4395) );
  INVX1 U5818 ( .A(n4573), .Y(n4396) );
  INVX1 U5819 ( .A(n4573), .Y(n4397) );
  INVX1 U5820 ( .A(n4573), .Y(n4398) );
  INVX1 U5821 ( .A(n4573), .Y(n4399) );
  INVX1 U5822 ( .A(n4572), .Y(n4400) );
  INVX1 U5823 ( .A(n4572), .Y(n4401) );
  INVX1 U5824 ( .A(n4572), .Y(n4402) );
  INVX1 U5825 ( .A(n4572), .Y(n4403) );
  INVX1 U5826 ( .A(n4572), .Y(n4404) );
  INVX1 U5827 ( .A(n4572), .Y(n4405) );
  INVX1 U5828 ( .A(n4572), .Y(n4406) );
  INVX1 U5829 ( .A(n4572), .Y(n4407) );
  INVX1 U5830 ( .A(n4572), .Y(n4408) );
  INVX1 U5831 ( .A(n4572), .Y(n4409) );
  INVX1 U5832 ( .A(n4571), .Y(n4410) );
  INVX1 U5833 ( .A(n4571), .Y(n4411) );
  INVX1 U5834 ( .A(n4571), .Y(n4412) );
  INVX1 U5835 ( .A(n4571), .Y(n4413) );
  INVX1 U5836 ( .A(n4571), .Y(n4414) );
  INVX1 U5837 ( .A(n4571), .Y(n4415) );
  INVX1 U5838 ( .A(n4571), .Y(n4416) );
  INVX1 U5839 ( .A(n4571), .Y(n4417) );
  INVX1 U5840 ( .A(n4570), .Y(n4418) );
  INVX1 U5841 ( .A(n4570), .Y(n4419) );
  INVX1 U5842 ( .A(n4570), .Y(n4420) );
  INVX1 U5843 ( .A(n4570), .Y(n4421) );
  INVX1 U5844 ( .A(n4570), .Y(n4422) );
  INVX1 U5845 ( .A(n4570), .Y(n4423) );
  INVX1 U5846 ( .A(n4570), .Y(n4424) );
  INVX1 U5847 ( .A(n4569), .Y(n4425) );
  INVX1 U5848 ( .A(n4570), .Y(n4426) );
  INVX1 U5849 ( .A(n4569), .Y(n4427) );
  INVX1 U5850 ( .A(n4569), .Y(n4428) );
  INVX1 U5851 ( .A(n4569), .Y(n4429) );
  INVX1 U5852 ( .A(n4569), .Y(n4430) );
  INVX1 U5853 ( .A(n4569), .Y(n4431) );
  INVX1 U5854 ( .A(n4569), .Y(n4432) );
  INVX1 U5855 ( .A(n4569), .Y(n4433) );
  INVX1 U5856 ( .A(n4568), .Y(n4434) );
  INVX1 U5857 ( .A(n4568), .Y(n4435) );
  INVX1 U5858 ( .A(n4568), .Y(n4436) );
  INVX1 U5859 ( .A(n4568), .Y(n4437) );
  INVX1 U5860 ( .A(n4568), .Y(n4438) );
  INVX1 U5861 ( .A(n4568), .Y(n4439) );
  INVX1 U5862 ( .A(n4568), .Y(n4440) );
  INVX1 U5863 ( .A(n4567), .Y(n4441) );
  INVX1 U5864 ( .A(n4568), .Y(n4442) );
  INVX1 U5865 ( .A(n4567), .Y(n4443) );
  INVX1 U5866 ( .A(n4567), .Y(n4444) );
  INVX1 U5867 ( .A(n4567), .Y(n4445) );
  INVX1 U5868 ( .A(n4567), .Y(n4446) );
  INVX1 U5869 ( .A(n4567), .Y(n4447) );
  INVX1 U5870 ( .A(n4567), .Y(n4448) );
  INVX1 U5871 ( .A(n4567), .Y(n4449) );
  INVX1 U5872 ( .A(n4567), .Y(n4450) );
  INVX1 U5873 ( .A(n4566), .Y(n4451) );
  INVX1 U5874 ( .A(n4567), .Y(n4452) );
  INVX1 U5875 ( .A(n4566), .Y(n4453) );
  INVX1 U5876 ( .A(n4566), .Y(n4454) );
  INVX1 U5877 ( .A(n4566), .Y(n4455) );
  INVX1 U5878 ( .A(n4566), .Y(n4456) );
  INVX1 U5879 ( .A(n4566), .Y(n4457) );
  INVX1 U5880 ( .A(n4566), .Y(n4458) );
  INVX1 U5881 ( .A(n4566), .Y(n4459) );
  INVX1 U5882 ( .A(n4566), .Y(n4460) );
  INVX1 U5883 ( .A(n4566), .Y(n4461) );
  INVX1 U5884 ( .A(n4565), .Y(n4462) );
  INVX1 U5885 ( .A(n4565), .Y(n4463) );
  INVX1 U5886 ( .A(n4565), .Y(n4464) );
  INVX1 U5887 ( .A(n4565), .Y(n4465) );
  INVX1 U5888 ( .A(n4565), .Y(n4466) );
  INVX1 U5889 ( .A(n4571), .Y(n4467) );
  INVX1 U5890 ( .A(n4579), .Y(n4468) );
  INVX1 U5891 ( .A(n4578), .Y(n4469) );
  INVX1 U5892 ( .A(n4578), .Y(n4470) );
  INVX1 U5893 ( .A(n4578), .Y(n4471) );
  INVX1 U5894 ( .A(n4570), .Y(n4472) );
  INVX1 U5895 ( .A(n4586), .Y(n4473) );
  INVX1 U5896 ( .A(n4578), .Y(n4474) );
  INVX1 U5897 ( .A(n4579), .Y(n4475) );
  INVX1 U5898 ( .A(n4581), .Y(n4476) );
  INVX1 U5899 ( .A(n4577), .Y(n4477) );
  INVX1 U5900 ( .A(n4583), .Y(n4478) );
  INVX1 U5901 ( .A(n4579), .Y(n4479) );
  INVX1 U5902 ( .A(n4584), .Y(n4480) );
  INVX1 U5903 ( .A(n4577), .Y(n4481) );
  INVX1 U5904 ( .A(n4569), .Y(n4482) );
  INVX1 U5905 ( .A(n4579), .Y(n4483) );
  INVX1 U5906 ( .A(n4581), .Y(n4484) );
  INVX1 U5907 ( .A(n4580), .Y(n4485) );
  INVX1 U5908 ( .A(n4585), .Y(n4486) );
  INVX1 U5909 ( .A(n4584), .Y(n4487) );
  INVX1 U5910 ( .A(n4585), .Y(n4488) );
  INVX1 U5911 ( .A(n4586), .Y(n4489) );
  INVX1 U5912 ( .A(n4584), .Y(n4490) );
  INVX1 U5913 ( .A(n4586), .Y(n4491) );
  INVX1 U5914 ( .A(n4580), .Y(n4492) );
  INVX1 U5915 ( .A(n4585), .Y(n4493) );
  INVX1 U5916 ( .A(n4584), .Y(n4494) );
  INVX1 U5917 ( .A(n4585), .Y(n4495) );
  INVX1 U5918 ( .A(n4584), .Y(n4496) );
  INVX1 U5919 ( .A(n4585), .Y(n4497) );
  INVX1 U5920 ( .A(n4584), .Y(n4498) );
  INVX1 U5921 ( .A(n4585), .Y(n4499) );
  INVX1 U5922 ( .A(n4579), .Y(n4500) );
  INVX1 U5923 ( .A(n4582), .Y(n4501) );
  INVX1 U5924 ( .A(n4577), .Y(n4502) );
  INVX1 U5925 ( .A(n4586), .Y(n4503) );
  INVX1 U5926 ( .A(n4577), .Y(n4504) );
  INVX1 U5927 ( .A(n4569), .Y(n4505) );
  INVX1 U5928 ( .A(n4577), .Y(n4506) );
  INVX1 U5929 ( .A(n4583), .Y(n4507) );
  INVX1 U5930 ( .A(n4584), .Y(n4508) );
  INVX1 U5931 ( .A(n4577), .Y(n4509) );
  INVX1 U5932 ( .A(n4568), .Y(n4510) );
  INVX1 U5933 ( .A(n4565), .Y(n4511) );
  INVX1 U5934 ( .A(n4580), .Y(n4512) );
  INVX1 U5935 ( .A(n4580), .Y(n4513) );
  INVX1 U5936 ( .A(n4583), .Y(n4514) );
  INVX1 U5937 ( .A(n4583), .Y(n4515) );
  INVX1 U5938 ( .A(n4583), .Y(n4516) );
  INVX1 U5939 ( .A(n4571), .Y(n4517) );
  INVX1 U5940 ( .A(n4580), .Y(n4518) );
  INVX1 U5941 ( .A(n4580), .Y(n4519) );
  INVX1 U5942 ( .A(n4577), .Y(n4520) );
  INVX1 U5943 ( .A(n4581), .Y(n4521) );
  INVX1 U5944 ( .A(n4581), .Y(n4522) );
  INVX1 U5945 ( .A(n4581), .Y(n4523) );
  INVX1 U5946 ( .A(n4586), .Y(n4524) );
  INVX1 U5947 ( .A(n4586), .Y(n4525) );
  INVX1 U5948 ( .A(n4586), .Y(n4526) );
  INVX1 U5949 ( .A(n4581), .Y(n4527) );
  INVX1 U5950 ( .A(n4581), .Y(n4528) );
  INVX1 U5951 ( .A(n4576), .Y(n4529) );
  INVX1 U5952 ( .A(n4576), .Y(n4530) );
  INVX1 U5953 ( .A(n4576), .Y(n4531) );
  INVX1 U5954 ( .A(n4576), .Y(n4532) );
  INVX1 U5955 ( .A(n4576), .Y(n4533) );
  INVX1 U5956 ( .A(n4576), .Y(n4534) );
  INVX1 U5957 ( .A(n4576), .Y(n4535) );
  INVX1 U5958 ( .A(n4576), .Y(n4536) );
  INVX1 U5959 ( .A(n4576), .Y(n4537) );
  INVX1 U5960 ( .A(n4576), .Y(n4538) );
  INVX1 U5961 ( .A(n4578), .Y(n4539) );
  INVX1 U5962 ( .A(n4579), .Y(n4540) );
  INVX1 U5963 ( .A(n4578), .Y(n4541) );
  INVX1 U5964 ( .A(n4579), .Y(n4542) );
  INVX1 U5965 ( .A(n4583), .Y(n4543) );
  INVX1 U5966 ( .A(n4583), .Y(n4544) );
  INVX1 U5967 ( .A(n4585), .Y(n4545) );
  INVX1 U5968 ( .A(n4580), .Y(n4546) );
  INVX1 U5969 ( .A(n4577), .Y(n4547) );
  INVX1 U5970 ( .A(n4578), .Y(n4548) );
  INVX1 U5971 ( .A(n4582), .Y(n4549) );
  INVX1 U5972 ( .A(n4582), .Y(n4550) );
  INVX1 U5973 ( .A(n4582), .Y(n4551) );
  INVX1 U5974 ( .A(n4582), .Y(n4552) );
  INVX1 U5975 ( .A(n4582), .Y(n4553) );
  INVX1 U5976 ( .A(n4582), .Y(n4554) );
  INVX1 U5977 ( .A(n4578), .Y(n4555) );
  INVX1 U5978 ( .A(n4582), .Y(n4556) );
  INVX1 U5979 ( .A(n4570), .Y(n4557) );
  INVX1 U5980 ( .A(n4579), .Y(n4558) );
  INVX1 U5981 ( .A(n4580), .Y(n4559) );
  INVX1 U5982 ( .A(n4577), .Y(n4560) );
  INVX1 U5983 ( .A(n4583), .Y(n4561) );
  INVX1 U5984 ( .A(n4568), .Y(n4562) );
  INVX1 U5985 ( .A(n4586), .Y(n4563) );
  INVX1 U5986 ( .A(n4565), .Y(n4564) );
endmodule


module aes_sbox ( sboxw, new_sboxw );
  input [31:0] sboxw;
  output [31:0] new_sboxw;
  wire   n1676, n1677, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n254, n255,
         n256, n257, n258, n259, n261, n262, n263, n264, n265, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n253, n260, n266, n352, n374, n929, n1345, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675;

  BUFX2 U1 ( .A(sboxw[11]), .Y(n102) );
  NAND2X1 U2 ( .A(sboxw[9]), .B(n51), .Y(n238) );
  INVX1 U3 ( .A(sboxw[9]), .Y(n207) );
  BUFX2 U4 ( .A(n261), .Y(n137) );
  OAI22XL U5 ( .A0(n136), .A1(n259), .B0(n1435), .B1(n141), .Y(n1434) );
  NAND2X1 U6 ( .A(n1562), .B(n100), .Y(n251) );
  BUFX2 U7 ( .A(n251), .Y(n138) );
  INVX1 U8 ( .A(n134), .Y(n135) );
  OAI21XL U9 ( .A0(n1439), .A1(n1440), .B0(sboxw[13]), .Y(n1438) );
  OAI221XL U10 ( .A0(n1585), .A1(n1289), .B0(n1587), .B1(n283), .C0(n254), .Y(
        n1439) );
  OAI222XL U11 ( .A0(n50), .A1(n239), .B0(sboxw[13]), .B1(n1431), .C0(n1432), 
        .C1(n169), .Y(n1427) );
  OAI222XL U12 ( .A0(n791), .A1(n566), .B0(n792), .B1(n568), .C0(sboxw[31]), 
        .C1(n793), .Y(new_sboxw[27]) );
  OAI222XL U13 ( .A0(n823), .A1(n566), .B0(n824), .B1(n568), .C0(sboxw[31]), 
        .C1(n825), .Y(new_sboxw[26]) );
  OAI222XL U14 ( .A0(n715), .A1(n568), .B0(sboxw[31]), .B1(n716), .C0(n717), 
        .C1(n566), .Y(new_sboxw[29]) );
  OAI222XL U15 ( .A0(n565), .A1(n566), .B0(n567), .B1(n568), .C0(sboxw[31]), 
        .C1(n569), .Y(new_sboxw[31]) );
  INVX1 U16 ( .A(sboxw[8]), .Y(n96) );
  INVX1 U17 ( .A(n96), .Y(n97) );
  AND2X2 U18 ( .A(n935), .B(n144), .Y(n1) );
  INVX1 U19 ( .A(n103), .Y(n1568) );
  NAND2X1 U20 ( .A(n101), .B(n44), .Y(n284) );
  BUFX12 U21 ( .A(n1676), .Y(new_sboxw[6]) );
  OAI2BB2XL U22 ( .B0(sboxw[7]), .B1(n404), .A0N(sboxw[7]), .A1N(n405), .Y(
        n1676) );
  BUFX12 U23 ( .A(n1677), .Y(new_sboxw[0]) );
  OAI2BB2XL U24 ( .B0(n1468), .B1(n1588), .A0N(n1469), .A1N(n1588), .Y(n1677)
         );
  OAI211X1 U25 ( .A0(n1411), .A1(n1266), .B0(n1412), .C0(n1413), .Y(
        new_sboxw[11]) );
  NAND2X1 U26 ( .A(n1580), .B(n99), .Y(n252) );
  NAND2XL U27 ( .A(n1583), .B(n45), .Y(n1326) );
  INVX1 U28 ( .A(n139), .Y(n1574) );
  INVX1 U29 ( .A(n207), .Y(n203) );
  NAND2XL U30 ( .A(n43), .B(n141), .Y(n317) );
  NAND2XL U31 ( .A(n1587), .B(n1558), .Y(n1339) );
  NAND2XL U32 ( .A(n48), .B(n1560), .Y(n1281) );
  INVXL U33 ( .A(n134), .Y(n136) );
  INVXL U34 ( .A(n288), .Y(n44) );
  NAND2XL U35 ( .A(n43), .B(n191), .Y(n254) );
  NAND2XL U36 ( .A(n138), .B(n139), .Y(n1359) );
  NAND2XL U37 ( .A(n1573), .B(n135), .Y(n1293) );
  NAND2XL U38 ( .A(n1553), .B(n1562), .Y(n269) );
  NAND2XL U39 ( .A(n1573), .B(n134), .Y(n1389) );
  NAND2XL U40 ( .A(n43), .B(n51), .Y(n246) );
  NAND2XL U41 ( .A(n1587), .B(n46), .Y(n1356) );
  NAND2XL U42 ( .A(n1560), .B(n169), .Y(n245) );
  NAND2X1 U43 ( .A(n77), .B(n179), .Y(n602) );
  NAND2X1 U44 ( .A(n34), .B(n164), .Y(n953) );
  INVX1 U45 ( .A(n89), .Y(n64) );
  AOI211XL U46 ( .A0(n1560), .A1(n141), .B0(n1461), .C0(n1307), .Y(n1460) );
  NAND2XL U47 ( .A(n337), .B(n135), .Y(n336) );
  AOI211XL U48 ( .A0(n1585), .A1(n1566), .B0(n307), .C0(n257), .Y(n1301) );
  NAND2XL U49 ( .A(n134), .B(n1566), .Y(n272) );
  NAND2XL U50 ( .A(n1562), .B(n1321), .Y(n1348) );
  AO22XL U51 ( .A0(n1582), .A1(n140), .B0(n1342), .B1(n1580), .Y(n1344) );
  NOR2XL U52 ( .A(n275), .B(n287), .Y(n240) );
  OAI21XL U53 ( .A0(n213), .A1(n951), .B0(n973), .Y(n1032) );
  INVX1 U54 ( .A(sboxw[26]), .Y(n77) );
  INVX1 U55 ( .A(n109), .Y(n34) );
  AOI211XL U56 ( .A0(n1564), .A1(sboxw[9]), .B0(n1433), .C0(n1434), .Y(n1432)
         );
  NOR2XL U57 ( .A(n45), .B(n101), .Y(n326) );
  NAND2BXL U58 ( .AN(n287), .B(n101), .Y(n243) );
  NAND2X1 U59 ( .A(n205), .B(n52), .Y(n10) );
  NAND2XL U60 ( .A(n101), .B(n45), .Y(n305) );
  NAND2X1 U61 ( .A(n98), .B(n203), .Y(n4) );
  NAND2X1 U62 ( .A(n205), .B(n52), .Y(n5) );
  NOR4XL U63 ( .A(n1328), .B(n1329), .C(n1574), .D(n1292), .Y(n1312) );
  AOI211XL U64 ( .A0(n48), .A1(n1566), .B0(n1572), .C0(n1575), .Y(n276) );
  OAI22XL U65 ( .A0(n287), .A1(n238), .B0(n203), .B1(n284), .Y(n328) );
  AO21XL U66 ( .A0(n43), .A1(n204), .B0(n1283), .Y(n1280) );
  NOR2XL U67 ( .A(n138), .B(n205), .Y(n1292) );
  AOI2BB2XL U68 ( .B0(n205), .B1(n1573), .A0N(n138), .A1N(n141), .Y(n1308) );
  AOI2BB1XL U69 ( .A0N(n170), .A1N(n288), .B0(n1298), .Y(n1393) );
  NAND2X1 U70 ( .A(n111), .B(n1534), .Y(n1071) );
  INVX1 U71 ( .A(n215), .Y(n213) );
  AOI2BB1X1 U72 ( .A0N(n265), .A1N(n14), .B0(n227), .Y(n264) );
  INVX1 U73 ( .A(n220), .Y(n218) );
  INVX1 U74 ( .A(n210), .Y(n208) );
  INVX1 U75 ( .A(n260), .Y(n223) );
  INVX1 U76 ( .A(n110), .Y(n1534) );
  AO22XL U77 ( .A0(n1580), .A1(n97), .B0(n5), .B1(n44), .Y(n286) );
  AO21XL U78 ( .A0(n205), .A1(n1560), .B0(n257), .Y(n1343) );
  OAI211XL U79 ( .A0(n251), .A1(n267), .B0(n272), .C0(n273), .Y(n271) );
  OAI22XL U80 ( .A0(n116), .A1(n218), .B0(n77), .B1(n158), .Y(n682) );
  OAI22XL U81 ( .A0(n108), .A1(n208), .B0(n34), .B1(n147), .Y(n1033) );
  OAI22XL U82 ( .A0(n266), .A1(n115), .B0(n117), .B1(n574), .Y(n674) );
  OAI22XL U83 ( .A0(n216), .A1(n107), .B0(n109), .B1(n147), .Y(n1025) );
  NOR2XL U84 ( .A(n137), .B(n203), .Y(n1298) );
  AOI21XL U85 ( .A0(n206), .A1(n1580), .B0(n1579), .Y(n285) );
  NAND2X1 U86 ( .A(n119), .B(n1668), .Y(n752) );
  NAND2X1 U87 ( .A(n121), .B(n77), .Y(n747) );
  NAND2X1 U88 ( .A(n113), .B(n34), .Y(n1066) );
  INVX1 U89 ( .A(n118), .Y(n1668) );
  INVX1 U90 ( .A(n99), .Y(n100) );
  INVX1 U91 ( .A(n88), .Y(n90) );
  NAND2XL U92 ( .A(n97), .B(n207), .Y(n334) );
  INVX1 U93 ( .A(n88), .Y(n89) );
  OAI222XL U94 ( .A0(n916), .A1(n917), .B0(n918), .B1(n919), .C0(sboxw[23]), 
        .C1(n920), .Y(new_sboxw[23]) );
  NOR4BXL U95 ( .AN(n254), .B(n255), .C(n256), .D(n257), .Y(n226) );
  NAND4BXL U96 ( .AN(n1362), .B(n254), .C(n302), .D(n1363), .Y(n1361) );
  OAI22XL U97 ( .A0(sboxw[31]), .A1(n754), .B0(n755), .B1(n1631), .Y(
        new_sboxw[28]) );
  OAI2BB2XL U98 ( .B0(n885), .B1(n1631), .A0N(n886), .A1N(n1631), .Y(
        new_sboxw[24]) );
  OAI2BB2XL U99 ( .B0(sboxw[31]), .B1(n630), .A0N(sboxw[31]), .A1N(n631), .Y(
        new_sboxw[30]) );
  OAI2BB2XL U100 ( .B0(n855), .B1(n1631), .A0N(n856), .A1N(n1631), .Y(
        new_sboxw[25]) );
  INVX1 U101 ( .A(n115), .Y(n116) );
  INVX1 U102 ( .A(n107), .Y(n108) );
  INVX1 U103 ( .A(n115), .Y(n117) );
  INVX1 U104 ( .A(n107), .Y(n109) );
  INVX1 U105 ( .A(sboxw[2]), .Y(n88) );
  INVX1 U106 ( .A(sboxw[10]), .Y(n99) );
  INVX1 U107 ( .A(sboxw[1]), .Y(n202) );
  INVX1 U108 ( .A(sboxw[26]), .Y(n115) );
  INVX1 U109 ( .A(sboxw[18]), .Y(n107) );
  INVX1 U110 ( .A(n504), .Y(n1618) );
  NAND2X1 U111 ( .A(n1652), .B(n185), .Y(n653) );
  NAND2X1 U112 ( .A(n1518), .B(n181), .Y(n1004) );
  NAND2X1 U113 ( .A(n1660), .B(n1642), .Y(n623) );
  BUFX2 U114 ( .A(n1587), .Y(n172) );
  NAND2X1 U115 ( .A(n1504), .B(n40), .Y(n974) );
  BUFX2 U116 ( .A(n13), .Y(n50) );
  NOR2X1 U117 ( .A(n1574), .B(n43), .Y(n1435) );
  INVX1 U118 ( .A(n322), .Y(n1550) );
  INVX1 U119 ( .A(n15), .Y(n21) );
  NAND2X1 U120 ( .A(n1604), .B(n176), .Y(n445) );
  BUFX2 U121 ( .A(n175), .Y(n176) );
  INVX1 U122 ( .A(n132), .Y(n1609) );
  BUFX2 U123 ( .A(n1620), .Y(n62) );
  NAND2X1 U124 ( .A(n176), .B(n59), .Y(n504) );
  NAND2X1 U125 ( .A(n56), .B(n1596), .Y(n381) );
  OAI22XL U126 ( .A0(n21), .A1(n349), .B0(n66), .B1(n403), .Y(n563) );
  OAI21XL U127 ( .A0(n178), .A1(n629), .B0(n671), .Y(n832) );
  OAI21XL U128 ( .A0(n167), .A1(n980), .B0(n1022), .Y(n1181) );
  BUFX2 U129 ( .A(n177), .Y(n178) );
  BUFX2 U130 ( .A(n166), .Y(n167) );
  INVX1 U131 ( .A(n188), .Y(n185) );
  INVX1 U132 ( .A(n1), .Y(n181) );
  NAND2X1 U133 ( .A(n1616), .B(n69), .Y(n530) );
  NAND2X1 U134 ( .A(n1656), .B(n178), .Y(n671) );
  NAND2X1 U135 ( .A(n1513), .B(n167), .Y(n1022) );
  NAND2X1 U136 ( .A(n1564), .B(n13), .Y(n327) );
  NAND2X1 U137 ( .A(n83), .B(n1661), .Y(n607) );
  BUFX2 U138 ( .A(n188), .Y(n187) );
  BUFX2 U139 ( .A(n1642), .Y(n72) );
  INVX1 U140 ( .A(n762), .Y(n1635) );
  INVX1 U141 ( .A(n1081), .Y(n1528) );
  INVX1 U142 ( .A(n464), .Y(n1615) );
  BUFX2 U143 ( .A(n1642), .Y(n73) );
  BUFX2 U144 ( .A(n1541), .Y(n39) );
  BUFX2 U145 ( .A(n1541), .Y(n40) );
  NAND2X1 U146 ( .A(n1595), .B(n1629), .Y(n397) );
  BUFX2 U147 ( .A(n1651), .Y(n76) );
  BUFX2 U148 ( .A(n1529), .Y(n33) );
  INVX1 U149 ( .A(n783), .Y(n1636) );
  INVX1 U150 ( .A(n1102), .Y(n1530) );
  INVX1 U151 ( .A(n163), .Y(n1652) );
  INVX1 U152 ( .A(n152), .Y(n1518) );
  INVX1 U153 ( .A(n188), .Y(n186) );
  INVX1 U154 ( .A(n184), .Y(n182) );
  INVX1 U155 ( .A(n901), .Y(n1660) );
  INVX1 U156 ( .A(n722), .Y(n1632) );
  INVX1 U157 ( .A(n1041), .Y(n1525) );
  INVX1 U158 ( .A(n743), .Y(n1634) );
  INVX1 U159 ( .A(n1062), .Y(n1521) );
  INVX1 U160 ( .A(n184), .Y(n183) );
  BUFX2 U161 ( .A(n1), .Y(n184) );
  NAND2X1 U162 ( .A(n1654), .B(n73), .Y(n788) );
  NAND2X1 U163 ( .A(n1526), .B(n39), .Y(n1107) );
  NAND2X1 U164 ( .A(n26), .B(n1505), .Y(n958) );
  INVX1 U165 ( .A(n822), .Y(n1643) );
  INVX1 U166 ( .A(n1171), .Y(n1520) );
  INVX1 U167 ( .A(n1250), .Y(n1504) );
  BUFX2 U168 ( .A(n44), .Y(n12) );
  NAND2X1 U169 ( .A(n6), .B(n1580), .Y(n322) );
  INVX1 U170 ( .A(n284), .Y(n43) );
  NOR2X1 U171 ( .A(n1560), .B(n1570), .Y(n1289) );
  NAND2X1 U172 ( .A(n189), .B(n1570), .Y(n1408) );
  BUFX2 U173 ( .A(n252), .Y(n139) );
  INVX1 U174 ( .A(n135), .Y(n1587) );
  NAND2X1 U175 ( .A(n1550), .B(n189), .Y(n1306) );
  INVX1 U176 ( .A(n316), .Y(n1564) );
  OAI21XL U177 ( .A0(n66), .A1(n423), .B0(n427), .Y(n1490) );
  INVX1 U178 ( .A(n402), .Y(n1604) );
  INVX1 U179 ( .A(n23), .Y(n24) );
  BUFX2 U180 ( .A(n1628), .Y(n67) );
  NAND2X1 U181 ( .A(n1609), .B(n23), .Y(n427) );
  INVX1 U182 ( .A(n431), .Y(n59) );
  BUFX2 U183 ( .A(n349), .Y(n132) );
  INVX1 U184 ( .A(n369), .Y(n1614) );
  INVX1 U185 ( .A(n482), .Y(n1608) );
  BUFX2 U186 ( .A(n1629), .Y(n68) );
  INVX1 U187 ( .A(n463), .Y(n55) );
  BUFX2 U188 ( .A(n1628), .Y(n66) );
  BUFX2 U189 ( .A(n1630), .Y(n175) );
  INVX1 U190 ( .A(n403), .Y(n1620) );
  INVX1 U191 ( .A(n376), .Y(n1596) );
  INVX1 U192 ( .A(n463), .Y(n56) );
  INVX1 U193 ( .A(n423), .Y(n1616) );
  BUFX2 U194 ( .A(n1629), .Y(n69) );
  INVX1 U195 ( .A(n1356), .Y(n1569) );
  INVX1 U196 ( .A(n1484), .Y(n1595) );
  INVX1 U197 ( .A(n711), .Y(n1599) );
  INVX1 U198 ( .A(n420), .Y(n1598) );
  NAND2X1 U199 ( .A(n176), .B(n60), .Y(n464) );
  OAI21XL U200 ( .A0(n70), .A1(n649), .B0(n653), .Y(n907) );
  OAI21XL U201 ( .A0(n38), .A1(n1000), .B0(n1004), .Y(n1256) );
  NAND2X1 U202 ( .A(n178), .B(n78), .Y(n762) );
  NAND2X1 U203 ( .A(n167), .B(n29), .Y(n1081) );
  OAI22XL U204 ( .A0(n187), .A1(n607), .B0(n608), .B1(n180), .Y(n606) );
  AOI211X1 U205 ( .A0(n1669), .A1(n154), .B0(n1636), .C0(n1638), .Y(n608) );
  INVX1 U206 ( .A(n588), .Y(n1638) );
  NAND2X1 U207 ( .A(n178), .B(n1663), .Y(n743) );
  NAND2X1 U208 ( .A(n167), .B(n1522), .Y(n1062) );
  NAND2X1 U209 ( .A(n178), .B(n1664), .Y(n783) );
  NAND2X1 U210 ( .A(n167), .B(n1531), .Y(n1102) );
  NAND2X1 U211 ( .A(n1663), .B(n154), .Y(n822) );
  NAND2X1 U212 ( .A(n1522), .B(n143), .Y(n1171) );
  NAND2X1 U213 ( .A(n178), .B(n80), .Y(n722) );
  NAND2X1 U214 ( .A(n167), .B(n31), .Y(n1041) );
  NAND2X1 U215 ( .A(n1661), .B(n1670), .Y(n901) );
  INVX1 U216 ( .A(n602), .Y(n1661) );
  INVX1 U217 ( .A(n953), .Y(n1505) );
  NAND2X1 U218 ( .A(n1662), .B(n74), .Y(n597) );
  NAND2X1 U219 ( .A(n1514), .B(n35), .Y(n948) );
  INVX1 U220 ( .A(n649), .Y(n1654) );
  INVX1 U221 ( .A(n1000), .Y(n1526) );
  NAND2X1 U222 ( .A(n6), .B(n12), .Y(n297) );
  INVX1 U223 ( .A(n628), .Y(n1656) );
  INVX1 U224 ( .A(n979), .Y(n1513) );
  INVX1 U225 ( .A(n1389), .Y(n1572) );
  NAND2X1 U226 ( .A(n1663), .B(n187), .Y(n679) );
  NAND2X1 U227 ( .A(n1522), .B(n184), .Y(n1030) );
  BUFX2 U228 ( .A(n575), .Y(n163) );
  BUFX2 U229 ( .A(n926), .Y(n152) );
  NAND2X1 U230 ( .A(n78), .B(n185), .Y(n736) );
  NAND2X1 U231 ( .A(n29), .B(n181), .Y(n1055) );
  INVX1 U232 ( .A(n311), .Y(n1548) );
  BUFX2 U233 ( .A(n1639), .Y(n71) );
  BUFX2 U234 ( .A(n1540), .Y(n38) );
  NAND2X1 U235 ( .A(n1581), .B(n49), .Y(n1357) );
  BUFX2 U236 ( .A(n1639), .Y(n70) );
  BUFX2 U237 ( .A(n1540), .Y(n37) );
  NOR2X1 U238 ( .A(n1662), .B(n1654), .Y(n573) );
  NOR2X1 U239 ( .A(n1514), .B(n1526), .Y(n924) );
  NOR2X1 U240 ( .A(n1605), .B(n1616), .Y(n347) );
  INVX1 U241 ( .A(n302), .Y(n1575) );
  INVX1 U242 ( .A(n721), .Y(n82) );
  INVX1 U243 ( .A(n1040), .Y(n26) );
  BUFX2 U244 ( .A(n1637), .Y(n177) );
  BUFX2 U245 ( .A(n1542), .Y(n166) );
  INVX1 U246 ( .A(n158), .Y(n74) );
  INVX1 U247 ( .A(n147), .Y(n35) );
  INVX1 U248 ( .A(n153), .Y(n1642) );
  INVX1 U249 ( .A(n935), .Y(n1541) );
  INVX1 U250 ( .A(n721), .Y(n83) );
  INVX1 U251 ( .A(n158), .Y(n75) );
  INVX1 U252 ( .A(n925), .Y(n36) );
  INVX1 U253 ( .A(n651), .Y(n1648) );
  INVX1 U254 ( .A(n1002), .Y(n1510) );
  INVX1 U255 ( .A(n629), .Y(n1651) );
  INVX1 U256 ( .A(n980), .Y(n1529) );
  INVX1 U257 ( .A(n844), .Y(n1647) );
  INVX1 U258 ( .A(n1193), .Y(n1503) );
  INVX1 U259 ( .A(n704), .Y(n1594) );
  INVX1 U260 ( .A(n1326), .Y(n1554) );
  INVX1 U261 ( .A(n241), .Y(n1552) );
  INVX1 U262 ( .A(n564), .Y(n1611) );
  INVX1 U263 ( .A(n868), .Y(n1653) );
  INVX1 U264 ( .A(n1217), .Y(n1519) );
  INVX1 U265 ( .A(n11), .Y(n525) );
  INVX1 U266 ( .A(n269), .Y(n1551) );
  INVX1 U267 ( .A(n646), .Y(n1657) );
  INVX1 U268 ( .A(n1123), .Y(n1610) );
  OAI22XL U269 ( .A0(n1), .A1(n958), .B0(n959), .B1(n1506), .Y(n957) );
  AOI211X1 U270 ( .A0(n1516), .A1(n143), .B0(n1530), .C0(n1527), .Y(n959) );
  INVX1 U271 ( .A(n939), .Y(n1527) );
  NOR3X1 U272 ( .A(n602), .B(n80), .C(n178), .Y(n843) );
  NOR3X1 U273 ( .A(n953), .B(n31), .C(n167), .Y(n1192) );
  NAND2X1 U274 ( .A(n1505), .B(n1533), .Y(n1250) );
  INVX1 U275 ( .A(n851), .Y(n1658) );
  INVX1 U276 ( .A(n1200), .Y(n1508) );
  INVX1 U277 ( .A(n997), .Y(n1507) );
  NOR2X1 U278 ( .A(n287), .B(n13), .Y(n330) );
  NAND2X1 U279 ( .A(n136), .B(n99), .Y(n303) );
  NAND3X1 U280 ( .A(n1334), .B(n104), .C(n12), .Y(n1430) );
  INVX1 U281 ( .A(n337), .Y(n1563) );
  INVX1 U282 ( .A(n267), .Y(n13) );
  INVX1 U283 ( .A(n249), .Y(n1570) );
  INVX1 U284 ( .A(n4), .Y(n189) );
  NAND2X1 U285 ( .A(n136), .B(n104), .Y(n1276) );
  INVX1 U286 ( .A(n1315), .Y(n1546) );
  NAND2X1 U287 ( .A(n99), .B(n45), .Y(n259) );
  INVX1 U288 ( .A(n137), .Y(n1562) );
  INVX1 U289 ( .A(n287), .Y(n1580) );
  BUFX2 U290 ( .A(n1585), .Y(n49) );
  INVX1 U291 ( .A(n1288), .Y(n1583) );
  INVX1 U292 ( .A(n138), .Y(n1560) );
  BUFX2 U293 ( .A(n104), .Y(n169) );
  BUFX2 U294 ( .A(n170), .Y(n171) );
  BUFX2 U295 ( .A(n1586), .Y(n170) );
  NAND2X1 U296 ( .A(n1493), .B(n128), .Y(n1478) );
  NAND2X1 U297 ( .A(n193), .B(n61), .Y(n369) );
  NAND2X1 U298 ( .A(n358), .B(n125), .Y(n23) );
  NAND2X1 U299 ( .A(n1607), .B(n63), .Y(n402) );
  NOR2X1 U300 ( .A(n21), .B(n19), .Y(n387) );
  NAND2X1 U301 ( .A(n55), .B(n63), .Y(n349) );
  OAI21XL U302 ( .A0(n176), .A1(n1608), .B0(n16), .Y(n1498) );
  NAND2X1 U303 ( .A(n127), .B(n64), .Y(n430) );
  NOR2X1 U304 ( .A(n127), .B(n396), .Y(n11) );
  NAND2X1 U305 ( .A(n60), .B(n64), .Y(n423) );
  NAND2X1 U306 ( .A(n64), .B(n1597), .Y(n376) );
  NAND2X1 U307 ( .A(n1613), .B(n15), .Y(n453) );
  NAND2X1 U308 ( .A(n8), .B(n64), .Y(n403) );
  NAND2X1 U309 ( .A(n430), .B(n16), .Y(n438) );
  NOR2X1 U310 ( .A(n24), .B(n396), .Y(n391) );
  INVX1 U311 ( .A(n494), .Y(n60) );
  NAND2X1 U312 ( .A(n1621), .B(n193), .Y(n443) );
  INVX1 U313 ( .A(n494), .Y(n61) );
  INVX1 U314 ( .A(n129), .Y(n1605) );
  INVX1 U315 ( .A(n419), .Y(n1607) );
  INVX1 U316 ( .A(n396), .Y(n1621) );
  INVX1 U317 ( .A(n358), .Y(n1629) );
  INVX1 U318 ( .A(n16), .Y(n1628) );
  INVX1 U319 ( .A(n441), .Y(n1630) );
  INVX1 U320 ( .A(n1492), .Y(n1602) );
  AOI221XL U321 ( .A0(n59), .A1(n65), .B0(n1478), .B1(n1607), .C0(n387), .Y(
        n1492) );
  OAI21XL U322 ( .A0(n125), .A1(n403), .B0(n453), .Y(n1483) );
  NOR2X1 U323 ( .A(n396), .B(n20), .Y(n472) );
  NAND2X1 U324 ( .A(n61), .B(n1600), .Y(n711) );
  OAI222XL U325 ( .A0(n18), .A1(n129), .B0(n69), .B1(n132), .C0(n1630), .C1(
        n131), .Y(n1482) );
  NAND2X1 U326 ( .A(n1607), .B(n1600), .Y(n420) );
  NAND2X1 U327 ( .A(n1596), .B(n8), .Y(n1484) );
  NAND2X1 U328 ( .A(n1601), .B(n174), .Y(n704) );
  NOR2X1 U329 ( .A(n16), .B(n463), .Y(n378) );
  NAND2X1 U330 ( .A(n66), .B(n63), .Y(n426) );
  INVX1 U331 ( .A(n425), .Y(n1601) );
  INVX1 U332 ( .A(n353), .Y(n1624) );
  OAI31XL U333 ( .A0(n1569), .A1(n1562), .A2(n278), .B0(n1553), .Y(n1367) );
  OAI211X1 U334 ( .A0(n193), .A1(n425), .B0(n426), .C0(n427), .Y(n421) );
  OAI21XL U335 ( .A0(n52), .A1(n282), .B0(n1293), .Y(n1291) );
  AOI222XL U336 ( .A0(n1609), .A1(n16), .B0(n1601), .B1(n66), .C0(n62), .C1(
        n65), .Y(n532) );
  NAND2X1 U337 ( .A(n1554), .B(n169), .Y(n311) );
  OAI22XL U338 ( .A0(n67), .A1(n711), .B0(n1120), .B1(n1597), .Y(n1117) );
  AOI2BB2X1 U339 ( .B0(n59), .B1(n194), .A0N(n131), .A1N(n69), .Y(n1120) );
  INVX1 U340 ( .A(n1293), .Y(n1571) );
  NOR2X1 U341 ( .A(n1579), .B(n1564), .Y(n250) );
  NAND2X1 U342 ( .A(n80), .B(n77), .Y(n649) );
  NAND2X1 U343 ( .A(n31), .B(n34), .Y(n1000) );
  OAI22XL U344 ( .A0(n249), .A1(n51), .B0(n170), .B1(n250), .Y(n248) );
  OAI21XL U345 ( .A0(n144), .A1(n980), .B0(n1030), .Y(n1249) );
  OAI22XL U346 ( .A0(n175), .A1(n130), .B0(n21), .B1(n402), .Y(n1138) );
  AOI211X1 U347 ( .A0(n1604), .A1(n1629), .B0(n466), .C0(n467), .Y(n465) );
  AOI2BB1X1 U348 ( .A0N(n1605), .A1N(n62), .B0(n127), .Y(n467) );
  NOR2X1 U349 ( .A(n162), .B(n185), .Y(n730) );
  NOR2X1 U350 ( .A(n151), .B(n181), .Y(n1049) );
  NAND2X1 U351 ( .A(n176), .B(n1613), .Y(n485) );
  NAND2X1 U352 ( .A(n1669), .B(n77), .Y(n628) );
  NAND2X1 U353 ( .A(n1516), .B(n34), .Y(n979) );
  OAI22XL U354 ( .A0(n101), .A1(n52), .B0(n189), .B1(n99), .Y(n306) );
  OAI22XL U355 ( .A0(n1637), .A1(n594), .B0(n185), .B1(n628), .Y(n883) );
  OAI22XL U356 ( .A0(n166), .A1(n945), .B0(n181), .B1(n979), .Y(n1232) );
  OAI22XL U357 ( .A0(n185), .A1(n753), .B0(n187), .B1(n628), .Y(n835) );
  OAI22XL U358 ( .A0(n181), .A1(n148), .B0(n184), .B1(n979), .Y(n1184) );
  INVX1 U359 ( .A(n909), .Y(n1640) );
  AOI221XL U360 ( .A0(n79), .A1(n74), .B0(n895), .B1(n1669), .C0(n613), .Y(
        n909) );
  INVX1 U361 ( .A(n1258), .Y(n1511) );
  AOI221XL U362 ( .A0(n30), .A1(n35), .B0(n1244), .B1(n1516), .C0(n964), .Y(
        n1258) );
  OAI21XL U363 ( .A0(n1558), .A1(n1573), .B0(n52), .Y(n1324) );
  NAND2X1 U364 ( .A(n1553), .B(n46), .Y(n241) );
  OAI21XL U365 ( .A0(n18), .A1(n126), .B0(n478), .Y(n476) );
  NAND2X1 U366 ( .A(n78), .B(n157), .Y(n588) );
  NAND2X1 U367 ( .A(n29), .B(n146), .Y(n939) );
  NOR2X1 U368 ( .A(n133), .B(n267), .Y(n257) );
  NOR2X1 U369 ( .A(n162), .B(n187), .Y(n617) );
  NOR2X1 U370 ( .A(n151), .B(n184), .Y(n968) );
  OAI222XL U371 ( .A0(n36), .A1(n1072), .B0(n39), .B1(n926), .C0(n166), .C1(
        n973), .Y(n1248) );
  OA21XL U372 ( .A0(n67), .A1(n130), .B0(n372), .Y(n401) );
  NAND4BX1 U373 ( .AN(n1576), .B(n1281), .C(n246), .D(n1389), .Y(n1395) );
  NAND2X1 U374 ( .A(n1669), .B(n1659), .Y(n646) );
  NAND2X1 U375 ( .A(n131), .B(n349), .Y(n1123) );
  NOR2X1 U376 ( .A(n185), .B(n600), .Y(n613) );
  NOR2X1 U377 ( .A(n181), .B(n150), .Y(n964) );
  OAI221XL U378 ( .A0(n190), .A1(n252), .B0(n1586), .B1(n133), .C0(n237), .Y(
        n1290) );
  NAND2X1 U379 ( .A(n1648), .B(n179), .Y(n844) );
  NAND2X1 U380 ( .A(n1510), .B(n164), .Y(n1193) );
  NAND2X1 U381 ( .A(n622), .B(n575), .Y(n868) );
  NAND2X1 U382 ( .A(n973), .B(n152), .Y(n1217) );
  NAND2X1 U383 ( .A(n1613), .B(n124), .Y(n564) );
  NAND2X1 U384 ( .A(n1649), .B(n87), .Y(n651) );
  NAND2X1 U385 ( .A(n1535), .B(n28), .Y(n1002) );
  OAI21XL U386 ( .A0(n21), .A1(n129), .B0(n401), .Y(n706) );
  NAND2X1 U387 ( .A(n441), .B(n174), .Y(n375) );
  INVX1 U388 ( .A(n329), .Y(n1556) );
  NAND2X1 U389 ( .A(n1579), .B(n267), .Y(n302) );
  NAND2X1 U390 ( .A(n82), .B(n115), .Y(n575) );
  NAND2X1 U391 ( .A(n26), .B(n107), .Y(n926) );
  NAND2X1 U392 ( .A(n1670), .B(n77), .Y(n629) );
  NAND2X1 U393 ( .A(n1533), .B(n34), .Y(n980) );
  OAI21XL U394 ( .A0(n178), .A1(n1667), .B0(n585), .Y(n915) );
  INVX1 U395 ( .A(n160), .Y(n1663) );
  INVX1 U396 ( .A(n149), .Y(n1522) );
  INVX1 U397 ( .A(n740), .Y(n1667) );
  INVX1 U398 ( .A(n1059), .Y(n1517) );
  NOR2X1 U399 ( .A(n51), .B(n137), .Y(n338) );
  NAND2X1 U400 ( .A(n1619), .B(n21), .Y(n478) );
  AOI2BB2X1 U401 ( .B0(n1263), .B1(n1506), .A0N(n147), .A1N(n979), .Y(n1262)
         );
  OAI221XL U402 ( .A0(n38), .A1(n1072), .B0(n1542), .B1(n945), .C0(n1090), .Y(
        n1263) );
  NOR2X1 U403 ( .A(n155), .B(n721), .Y(n604) );
  NOR2X1 U404 ( .A(n936), .B(n1040), .Y(n955) );
  NAND3X1 U405 ( .A(n438), .B(n174), .C(n55), .Y(n551) );
  NOR2X1 U406 ( .A(n128), .B(n130), .Y(n389) );
  INVX1 U407 ( .A(n162), .Y(n1664) );
  INVX1 U408 ( .A(n151), .Y(n1531) );
  INVX1 U409 ( .A(n753), .Y(n1662) );
  INVX1 U410 ( .A(n148), .Y(n1514) );
  OAI221XL U411 ( .A0(n71), .A1(n159), .B0(n1637), .B1(n594), .C0(n771), .Y(
        n914) );
  INVX1 U412 ( .A(n1040), .Y(n1523) );
  NAND2X1 U413 ( .A(n130), .B(n423), .Y(n1131) );
  INVX1 U414 ( .A(n283), .Y(n1558) );
  NOR2X1 U415 ( .A(n574), .B(n160), .Y(n615) );
  NOR2X1 U416 ( .A(n925), .B(n149), .Y(n966) );
  INVX1 U417 ( .A(n4), .Y(n190) );
  INVX1 U418 ( .A(n282), .Y(n1581) );
  INVX1 U419 ( .A(n156), .Y(n1669) );
  INVX1 U420 ( .A(n145), .Y(n1516) );
  NAND2X1 U421 ( .A(n1605), .B(n65), .Y(n371) );
  BUFX2 U422 ( .A(n584), .Y(n153) );
  INVX1 U423 ( .A(n752), .Y(n80) );
  INVX1 U424 ( .A(n1071), .Y(n31) );
  INVX1 U425 ( .A(n600), .Y(n1670) );
  INVX1 U426 ( .A(n150), .Y(n1533) );
  INVX1 U427 ( .A(n752), .Y(n81) );
  INVX1 U428 ( .A(n1071), .Y(n32) );
  BUFX2 U429 ( .A(n584), .Y(n154) );
  BUFX2 U430 ( .A(n935), .Y(n143) );
  INVX1 U431 ( .A(n579), .Y(n1649) );
  INVX1 U432 ( .A(n930), .Y(n1535) );
  INVX1 U433 ( .A(n657), .Y(n78) );
  INVX1 U434 ( .A(n1008), .Y(n29) );
  OAI222XL U435 ( .A0(n645), .A1(n155), .B0(n594), .B1(n153), .C0(n1644), .C1(
        n161), .Y(n642) );
  OAI222XL U436 ( .A0(n996), .A1(n936), .B0(n945), .B1(n142), .C0(n1539), .C1(
        n951), .Y(n993) );
  OA21XL U437 ( .A0(n45), .A1(n236), .B0(n245), .Y(n1277) );
  INVX1 U438 ( .A(n657), .Y(n79) );
  INVX1 U439 ( .A(n1008), .Y(n30) );
  INVX1 U440 ( .A(n155), .Y(n1639) );
  INVX1 U441 ( .A(n144), .Y(n1540) );
  BUFX2 U442 ( .A(n935), .Y(n142) );
  NAND2X1 U443 ( .A(n1605), .B(n174), .Y(n377) );
  OAI221XL U444 ( .A0(n187), .A1(n851), .B0(n186), .B1(n646), .C0(n612), .Y(
        n850) );
  OAI221XL U445 ( .A0(n1), .A1(n1200), .B0(n182), .B1(n997), .C0(n963), .Y(
        n1199) );
  BUFX2 U446 ( .A(n104), .Y(n168) );
  AOI32X1 U447 ( .A0(n482), .A1(n123), .A2(n1593), .B0(n1594), .B1(sboxw[0]), 
        .Y(n481) );
  OAI31XL U448 ( .A0(n1632), .A1(n1669), .A2(n1641), .B0(n1659), .Y(n732) );
  OAI31XL U449 ( .A0(n1525), .A1(n1516), .A2(n1537), .B0(n1509), .Y(n1051) );
  OAI211X1 U450 ( .A0(n578), .A1(n721), .B0(n722), .C0(n597), .Y(n719) );
  OAI211X1 U451 ( .A0(n183), .A1(n1040), .B0(n1041), .C0(n948), .Y(n1038) );
  OAI211X1 U452 ( .A0(n65), .A1(n347), .B0(n564), .C0(n525), .Y(n562) );
  BUFX2 U453 ( .A(n1585), .Y(n48) );
  INVX1 U454 ( .A(n667), .Y(n1637) );
  INVX1 U455 ( .A(n146), .Y(n1542) );
  INVX1 U456 ( .A(n578), .Y(n188) );
  NAND2X1 U457 ( .A(n153), .B(n585), .Y(n578) );
  INVX1 U458 ( .A(n272), .Y(n1565) );
  OAI2BB2XL U459 ( .B0(n645), .B1(n601), .A0N(n75), .A1N(n818), .Y(n817) );
  OAI2BB2XL U460 ( .B0(n996), .B1(n952), .A0N(n36), .A1N(n1167), .Y(n1166) );
  OAI21XL U461 ( .A0(n87), .A1(n602), .B0(n603), .Y(n599) );
  OAI21XL U462 ( .A0(n28), .A1(n953), .B0(n954), .Y(n950) );
  NAND2X1 U463 ( .A(n81), .B(n1659), .Y(n851) );
  NAND2X1 U464 ( .A(n32), .B(n1509), .Y(n1200) );
  NAND2X1 U465 ( .A(n1516), .B(n1509), .Y(n997) );
  NAND2X1 U466 ( .A(n157), .B(n77), .Y(n656) );
  NAND2X1 U467 ( .A(n146), .B(n34), .Y(n1007) );
  NAND2X1 U468 ( .A(n70), .B(n115), .Y(n652) );
  NAND2X1 U469 ( .A(n1540), .B(n107), .Y(n1003) );
  NAND2X1 U470 ( .A(n656), .B(n155), .Y(n664) );
  NAND2X1 U471 ( .A(n1007), .B(n936), .Y(n1015) );
  NAND3X1 U472 ( .A(n664), .B(n179), .C(n82), .Y(n809) );
  NAND3X1 U473 ( .A(n1015), .B(n164), .C(n26), .Y(n1158) );
  NOR2X1 U474 ( .A(n587), .B(n158), .Y(n724) );
  NOR2X1 U475 ( .A(n938), .B(n147), .Y(n1043) );
  NAND2X1 U476 ( .A(n667), .B(n179), .Y(n601) );
  NAND2X1 U477 ( .A(n146), .B(n164), .Y(n952) );
  NAND2X1 U478 ( .A(n818), .B(n157), .Y(n661) );
  NAND2X1 U479 ( .A(n1167), .B(n1018), .Y(n1012) );
  NAND2X1 U480 ( .A(n1662), .B(n179), .Y(n603) );
  NAND2X1 U481 ( .A(n1514), .B(n164), .Y(n954) );
  AO22X1 U482 ( .A0(n1675), .A1(n1632), .B0(n1661), .B1(n614), .Y(n620) );
  AO22X1 U483 ( .A0(n1506), .A1(n1525), .B0(n1505), .B1(n965), .Y(n971) );
  INVX1 U484 ( .A(n580), .Y(n1655) );
  INVX1 U485 ( .A(n931), .Y(n1512) );
  INVX1 U486 ( .A(n409), .Y(n1589) );
  INVX1 U487 ( .A(n595), .Y(n1646) );
  INVX1 U488 ( .A(n946), .Y(n1524) );
  NAND2X1 U489 ( .A(n169), .B(n41), .Y(n1315) );
  NAND2X1 U490 ( .A(n137), .B(n7), .Y(n337) );
  NAND2X1 U491 ( .A(n1582), .B(n1568), .Y(n288) );
  NAND2BX1 U492 ( .AN(n261), .B(n47), .Y(n283) );
  NOR2X1 U493 ( .A(n236), .B(n7), .Y(n1337) );
  NAND2X1 U494 ( .A(n140), .B(n238), .Y(n267) );
  NAND2X1 U495 ( .A(n9), .B(n99), .Y(n249) );
  INVX1 U496 ( .A(n103), .Y(n45) );
  NOR2X1 U497 ( .A(n1584), .B(n323), .Y(n1288) );
  INVX1 U498 ( .A(n238), .Y(n134) );
  AND2X2 U499 ( .A(n47), .B(n104), .Y(n6) );
  INVX1 U500 ( .A(n6), .Y(n236) );
  INVX1 U501 ( .A(n284), .Y(n1566) );
  NAND2X1 U502 ( .A(n12), .B(n47), .Y(n316) );
  NAND2X1 U503 ( .A(n303), .B(n5), .Y(n1334) );
  BUFX2 U504 ( .A(n96), .Y(n52) );
  INVX1 U505 ( .A(n295), .Y(n1549) );
  BUFX2 U506 ( .A(n243), .Y(n133) );
  NAND2X1 U507 ( .A(n326), .B(n189), .Y(n1388) );
  BUFX2 U508 ( .A(n96), .Y(n51) );
  INVX1 U509 ( .A(n244), .Y(n1573) );
  INVX1 U510 ( .A(n10), .Y(n1586) );
  INVX1 U511 ( .A(n243), .Y(n1579) );
  INVX1 U512 ( .A(n140), .Y(n1585) );
  OAI31XL U513 ( .A0(n295), .A1(n45), .A2(n51), .B0(n1430), .Y(n1429) );
  INVX1 U514 ( .A(n258), .Y(n1584) );
  BUFX2 U515 ( .A(n441), .Y(n127) );
  INVX1 U516 ( .A(n455), .Y(n1622) );
  NOR2BX1 U517 ( .AN(n453), .B(n454), .Y(n452) );
  OAI221XL U518 ( .A0(n67), .A1(n495), .B0(n176), .B1(n130), .C0(n513), .Y(
        n1497) );
  OAI211X1 U519 ( .A0(n1487), .A1(n173), .B0(n1488), .C0(n1484), .Y(n1486) );
  OAI221XL U520 ( .A0(n18), .A1(n402), .B0(n196), .B1(n129), .C0(n1491), .Y(
        n1489) );
  BUFX2 U521 ( .A(n368), .Y(n130) );
  NAND2X1 U522 ( .A(n126), .B(n494), .Y(n482) );
  NOR4BX1 U523 ( .AN(n355), .B(n428), .C(n429), .D(n62), .Y(n406) );
  OAI22XL U524 ( .A0(n16), .A1(n132), .B0(n56), .B1(n430), .Y(n429) );
  OAI222XL U525 ( .A0(n15), .A1(n130), .B0(n20), .B1(n431), .C0(n199), .C1(n19), .Y(n428) );
  BUFX2 U526 ( .A(n419), .Y(n126) );
  NAND2X1 U527 ( .A(n1623), .B(n57), .Y(n463) );
  BUFX2 U528 ( .A(n1597), .Y(n174) );
  BUFX2 U529 ( .A(n359), .Y(n16) );
  BUFX2 U530 ( .A(n358), .Y(n123) );
  INVX1 U531 ( .A(n431), .Y(n1619) );
  INVX1 U532 ( .A(n89), .Y(n63) );
  BUFX2 U533 ( .A(n348), .Y(n128) );
  BUFX2 U534 ( .A(n495), .Y(n129) );
  INVX1 U535 ( .A(n368), .Y(n1613) );
  INVX1 U536 ( .A(n197), .Y(n193) );
  BUFX2 U537 ( .A(n359), .Y(n125) );
  BUFX2 U538 ( .A(n396), .Y(n131) );
  INVX1 U539 ( .A(n700), .Y(n1626) );
  INVX1 U540 ( .A(n22), .Y(n448) );
  NAND2X1 U541 ( .A(n1621), .B(n195), .Y(n372) );
  NOR2X1 U542 ( .A(n529), .B(n1625), .Y(n353) );
  OAI22XL U543 ( .A0(n176), .A1(n129), .B0(n128), .B1(n442), .Y(n415) );
  NOR2X1 U544 ( .A(n19), .B(n489), .Y(n411) );
  NAND2X1 U545 ( .A(n174), .B(n53), .Y(n409) );
  INVX1 U546 ( .A(n512), .Y(n1625) );
  NAND2X1 U547 ( .A(n1624), .B(n58), .Y(n425) );
  INVX1 U548 ( .A(n489), .Y(n1600) );
  INVX1 U549 ( .A(n348), .Y(n65) );
  BUFX2 U550 ( .A(n1597), .Y(n173) );
  AOI222XL U551 ( .A0(n344), .A1(n54), .B0(n1592), .B1(n345), .C0(n1591), .C1(
        n346), .Y(n343) );
  NAND4X1 U552 ( .A(n355), .B(n132), .C(n356), .D(n357), .Y(n345) );
  NAND4BX1 U553 ( .AN(n363), .B(n364), .C(n365), .D(n366), .Y(n344) );
  OAI221XL U554 ( .A0(n347), .A1(n196), .B0(n348), .B1(n349), .C0(n350), .Y(
        n346) );
  INVX1 U555 ( .A(n196), .Y(n194) );
  AOI211X1 U556 ( .A0(n1595), .A1(n20), .B0(n1479), .C0(n1480), .Y(n1470) );
  OAI31XL U557 ( .A0(n398), .A1(n1608), .A2(n20), .B0(n701), .Y(n1480) );
  OAI222XL U558 ( .A0(n65), .A1(n381), .B0(n66), .B1(n704), .C0(n1481), .C1(
        n173), .Y(n1479) );
  NOR4X1 U559 ( .A(n1482), .B(n1483), .C(n1618), .D(n712), .Y(n1481) );
  INVX1 U560 ( .A(n398), .Y(n1593) );
  OAI22XL U561 ( .A0(n360), .A1(n463), .B0(n526), .B1(n376), .Y(n1119) );
  AOI221XL U562 ( .A0(n62), .A1(n123), .B0(n1621), .B1(n16), .C0(n360), .Y(
        n357) );
  OAI22XL U563 ( .A0(n10), .A1(n316), .B0(n44), .B1(n303), .Y(n1329) );
  OAI2BB2XL U564 ( .B0(n127), .B1(n552), .A0N(n441), .A1N(n411), .Y(n1118) );
  OAI2BB2XL U565 ( .B0(n136), .B1(n239), .A0N(n136), .A1N(n240), .Y(n233) );
  OAI222XL U566 ( .A0(n127), .A1(n495), .B0(n21), .B1(n403), .C0(n431), .C1(
        n359), .Y(n1121) );
  OAI222XL U567 ( .A0(n138), .A1(n136), .B0(n50), .B1(n139), .C0(n10), .C1(
        n244), .Y(n247) );
  OAI222XL U568 ( .A0(n244), .A1(n192), .B0(n249), .B1(n5), .C0(n13), .C1(n261), .Y(n255) );
  AOI222XL U569 ( .A0(n8), .A1(n456), .B0(n1604), .B1(n194), .C0(n59), .C1(n15), .Y(n547) );
  NAND4BX1 U570 ( .AN(n712), .B(n372), .C(n130), .D(n713), .Y(n709) );
  AOI222XL U571 ( .A0(n62), .A1(n15), .B0(n199), .B1(n714), .C0(n515), .C1(n18), .Y(n713) );
  NAND2X1 U572 ( .A(n463), .B(n442), .Y(n714) );
  NOR3X1 U573 ( .A(n489), .B(n68), .C(n463), .Y(n363) );
  OAI22XL U574 ( .A0(n195), .A1(n423), .B0(n67), .B1(n1610), .Y(n1122) );
  OAI222XL U575 ( .A0(n431), .A1(n123), .B0(n359), .B1(n423), .C0(n23), .C1(
        n126), .Y(n1124) );
  OAI22XL U576 ( .A0(n178), .A1(n753), .B0(n158), .B1(n668), .Y(n641) );
  OAI22XL U577 ( .A0(n167), .A1(n148), .B0(n147), .B1(n1019), .Y(n992) );
  OAI21XL U578 ( .A0(n223), .A1(n161), .B0(n622), .Y(n681) );
  AOI222XL U579 ( .A0(n67), .A1(n60), .B0(n529), .B1(n1630), .C0(n1604), .C1(
        n194), .Y(n528) );
  NAND2X1 U580 ( .A(n1668), .B(n86), .Y(n721) );
  NAND2X1 U581 ( .A(n1534), .B(n27), .Y(n1040) );
  OAI22XL U582 ( .A0(n134), .A1(n138), .B0(n140), .B1(n281), .Y(n1320) );
  OAI221XL U583 ( .A0(n24), .A1(n711), .B0(n23), .B1(n420), .C0(n386), .Y(n710) );
  OAI221XL U584 ( .A0(n141), .A1(n241), .B0(n50), .B1(n269), .C0(n1299), .Y(
        n1465) );
  AOI211X1 U585 ( .A0(n190), .A1(n46), .B0(n1455), .C0(n1456), .Y(n1450) );
  OAI22XL U586 ( .A0(n13), .A1(n251), .B0(n204), .B1(n139), .Y(n1456) );
  OAI221XL U587 ( .A0(n250), .A1(n334), .B0(n283), .B1(n267), .C0(n304), .Y(
        n1455) );
  NOR4BX1 U588 ( .AN(n1408), .B(n1452), .C(n1453), .D(n1572), .Y(n1451) );
  OAI21XL U589 ( .A0(n50), .A1(n316), .B0(n1339), .Y(n1453) );
  OAI221XL U590 ( .A0(n13), .A1(n283), .B0(n134), .B1(n284), .C0(n285), .Y(
        n279) );
  OAI22XL U591 ( .A0(n69), .A1(n423), .B0(n67), .B1(n512), .Y(n511) );
  OAI2BB2XL U592 ( .B0(n235), .B1(n236), .A0N(n237), .A1N(n12), .Y(n234) );
  OAI22XL U593 ( .A0(n189), .A1(n258), .B0(n51), .B1(n259), .Y(n256) );
  OAI22XL U594 ( .A0(n845), .A1(n179), .B0(n253), .B1(n810), .Y(n842) );
  AOI211X1 U595 ( .A0(n1654), .A1(n574), .B0(n846), .C0(n847), .Y(n845) );
  OAI21XL U596 ( .A0(n185), .A1(n753), .B0(n627), .Y(n846) );
  OAI31XL U597 ( .A0(n87), .A1(n73), .A2(n579), .B0(n671), .Y(n847) );
  OAI22XL U598 ( .A0(n1194), .A1(n164), .B0(n214), .B1(n1159), .Y(n1191) );
  AOI211X1 U599 ( .A0(n1526), .A1(n925), .B0(n1195), .C0(n1196), .Y(n1194) );
  OAI31XL U600 ( .A0(n28), .A1(n39), .A2(n930), .B0(n1022), .Y(n1196) );
  OAI21XL U601 ( .A0(n181), .A1(n148), .B0(n978), .Y(n1195) );
  NOR2X1 U602 ( .A(n787), .B(n1650), .Y(n579) );
  NOR2X1 U603 ( .A(n1106), .B(n1536), .Y(n930) );
  OAI22XL U604 ( .A0(n17), .A1(n128), .B0(n359), .B1(n442), .Y(n516) );
  OAI211X1 U605 ( .A0(n320), .A1(n169), .B0(n321), .C0(n322), .Y(n319) );
  NAND3X1 U606 ( .A(n172), .B(n1582), .C(n6), .Y(n321) );
  OAI22XL U607 ( .A0(n287), .A1(n334), .B0(n5), .B1(n281), .Y(n1397) );
  OAI22XL U608 ( .A0(n261), .A1(n10), .B0(n284), .B1(n192), .Y(n1323) );
  OAI22XL U609 ( .A0(n17), .A1(n195), .B0(n66), .B1(n463), .Y(n1139) );
  AOI222XL U610 ( .A0(n1574), .A1(n267), .B0(n204), .B1(n1467), .C0(n1555), 
        .C1(n49), .Y(n1466) );
  NAND2X1 U611 ( .A(n156), .B(n752), .Y(n740) );
  NAND2X1 U612 ( .A(n145), .B(n1071), .Y(n1059) );
  OAI22XL U613 ( .A0(n101), .A1(n49), .B0(n189), .B1(n47), .Y(n237) );
  NOR4X1 U614 ( .A(n728), .B(n729), .C(n730), .D(n1643), .Y(n727) );
  OAI2BB1X1 U615 ( .A0N(n1661), .A1N(n731), .B0(n607), .Y(n729) );
  OAI211X1 U616 ( .A0(n177), .A1(n575), .B0(n732), .C0(n733), .Y(n728) );
  OAI21XL U617 ( .A0(n74), .A1(n1668), .B0(n153), .Y(n731) );
  NOR4X1 U618 ( .A(n1047), .B(n1048), .C(n1049), .D(n1520), .Y(n1046) );
  OAI2BB1X1 U619 ( .A0N(n1505), .A1N(n1050), .B0(n958), .Y(n1048) );
  OAI211X1 U620 ( .A0(n166), .A1(n926), .B0(n1051), .C0(n1052), .Y(n1047) );
  OAI21XL U621 ( .A0(n35), .A1(n1534), .B0(n142), .Y(n1050) );
  AOI221XL U622 ( .A0(n65), .A1(n411), .B0(n1589), .B1(n517), .C0(n518), .Y(
        n496) );
  OAI22XL U623 ( .A0(n519), .A1(n54), .B0(n520), .B1(n407), .Y(n518) );
  NAND4X1 U624 ( .A(n530), .B(n372), .C(n531), .D(n532), .Y(n517) );
  AOI221XL U625 ( .A0(n1607), .A1(n20), .B0(n56), .B1(n124), .C0(n521), .Y(
        n520) );
  OAI22XL U626 ( .A0(n189), .A1(n249), .B0(n170), .B1(n258), .Y(n1396) );
  NAND2X1 U627 ( .A(n47), .B(n1582), .Y(n282) );
  OAI22XL U628 ( .A0(n161), .A1(n574), .B0(n585), .B1(n668), .Y(n774) );
  OAI22XL U629 ( .A0(n73), .A1(n649), .B0(n71), .B1(n770), .Y(n769) );
  OAI22XL U630 ( .A0(n39), .A1(n1000), .B0(n38), .B1(n1089), .Y(n1088) );
  OAI22XL U631 ( .A0(n973), .A1(n936), .B0(n208), .B1(n1072), .Y(n1150) );
  NOR4BX1 U632 ( .AN(n893), .B(n894), .C(n1663), .D(n730), .Y(n892) );
  OAI21XL U633 ( .A0(n1667), .A1(n656), .B0(n836), .Y(n894) );
  AOI222XL U634 ( .A0(n72), .A1(n76), .B0(n1637), .B1(n773), .C0(n219), .C1(
        n83), .Y(n893) );
  NOR4BX1 U635 ( .AN(n1242), .B(n1243), .C(n1522), .D(n1049), .Y(n1241) );
  OAI21XL U636 ( .A0(n1517), .A1(n1007), .B0(n1185), .Y(n1243) );
  AOI222XL U637 ( .A0(n40), .A1(n33), .B0(n1542), .B1(n1092), .C0(n209), .C1(
        n1523), .Y(n1242) );
  NOR4BX1 U638 ( .AN(n310), .B(n1458), .C(n1459), .D(n1548), .Y(n1442) );
  NOR3X1 U639 ( .A(n236), .B(n172), .C(n46), .Y(n1459) );
  OAI22XL U640 ( .A0(n1460), .A1(n104), .B0(n204), .B1(n239), .Y(n1458) );
  AOI2BB2X1 U641 ( .B0(n373), .B1(n124), .A0N(n19), .A1N(n375), .Y(n365) );
  NOR4BX1 U642 ( .AN(n701), .B(n702), .C(n703), .D(n1594), .Y(n684) );
  OAI22XL U643 ( .A0(n705), .A1(n174), .B0(n199), .B1(n552), .Y(n702) );
  AOI211X1 U644 ( .A0(n1616), .A1(n128), .B0(n706), .C0(n707), .Y(n705) );
  NOR4BX1 U645 ( .AN(n581), .B(n654), .C(n655), .D(n1651), .Y(n632) );
  OAI22XL U646 ( .A0(n155), .A1(n575), .B0(n83), .B1(n656), .Y(n655) );
  OAI222XL U647 ( .A0(n188), .A1(n594), .B0(n578), .B1(n657), .C0(n253), .C1(
        n161), .Y(n654) );
  NOR4BX1 U648 ( .AN(n932), .B(n1005), .C(n1006), .D(n1529), .Y(n983) );
  OAI22XL U649 ( .A0(n936), .A1(n926), .B0(n1523), .B1(n1007), .Y(n1006) );
  OAI222XL U650 ( .A0(n184), .A1(n945), .B0(n183), .B1(n1008), .C0(n214), .C1(
        n951), .Y(n1005) );
  NAND3X1 U651 ( .A(n359), .B(n57), .C(n353), .Y(n546) );
  OA21XL U652 ( .A0(n71), .A1(n160), .B0(n598), .Y(n627) );
  OA21XL U653 ( .A0(n38), .A1(n149), .B0(n949), .Y(n978) );
  NOR2X1 U654 ( .A(n52), .B(n7), .Y(n1283) );
  BUFX2 U655 ( .A(n1675), .Y(n179) );
  BUFX2 U656 ( .A(n165), .Y(n164) );
  BUFX2 U657 ( .A(n1506), .Y(n165) );
  NAND2X1 U658 ( .A(n1664), .B(n218), .Y(n669) );
  OAI222XL U659 ( .A0(n284), .A1(n267), .B0(n13), .B1(n244), .C0(n204), .C1(
        n287), .Y(n1328) );
  NAND2X1 U660 ( .A(n218), .B(n223), .Y(n584) );
  NAND2X1 U661 ( .A(n208), .B(n213), .Y(n935) );
  NOR3X1 U662 ( .A(n1283), .B(n330), .C(n1298), .Y(n1297) );
  NAND2BX1 U663 ( .AN(n431), .B(n441), .Y(n362) );
  AOI2BB2X1 U664 ( .B0(n199), .B1(n1613), .A0N(n1630), .A1N(n495), .Y(n693) );
  NAND2X1 U665 ( .A(n218), .B(n81), .Y(n595) );
  NAND2X1 U666 ( .A(n208), .B(n32), .Y(n946) );
  NAND2X1 U667 ( .A(n1656), .B(n223), .Y(n580) );
  NAND2X1 U668 ( .A(n1513), .B(n213), .Y(n931) );
  NAND4BX1 U669 ( .AN(n615), .B(n788), .C(n804), .D(n805), .Y(n794) );
  NAND3X1 U670 ( .A(n585), .B(n86), .C(n579), .Y(n804) );
  AOI222XL U671 ( .A0(n1670), .A1(n682), .B0(n1656), .B1(n219), .C0(n79), .C1(
        n187), .Y(n805) );
  NAND4BX1 U672 ( .AN(n966), .B(n1107), .C(n1153), .D(n1154), .Y(n1143) );
  NAND3X1 U673 ( .A(n144), .B(n27), .C(n930), .Y(n1153) );
  AOI222XL U674 ( .A0(n1533), .A1(n1033), .B0(n1513), .B1(n209), .C0(n30), 
        .C1(n1), .Y(n1154) );
  OA21XL U675 ( .A0(n196), .A1(n361), .B0(n362), .Y(n356) );
  NAND2X1 U676 ( .A(n1613), .B(n195), .Y(n514) );
  NAND4X1 U677 ( .A(n668), .B(n653), .C(n785), .D(n786), .Y(n780) );
  OAI2BB1X1 U678 ( .A0N(n650), .A1N(n161), .B0(n154), .Y(n785) );
  AOI222XL U679 ( .A0(n71), .A1(n80), .B0(n787), .B1(n177), .C0(n1656), .C1(
        n219), .Y(n786) );
  NAND4X1 U680 ( .A(n1019), .B(n1004), .C(n1104), .D(n1105), .Y(n1099) );
  OAI2BB1X1 U681 ( .A0N(n1001), .A1N(n951), .B0(n143), .Y(n1104) );
  AOI222XL U682 ( .A0(n38), .A1(n31), .B0(n1106), .B1(n166), .C0(n1513), .C1(
        n209), .Y(n1105) );
  OAI31XL U683 ( .A0(n389), .A1(n390), .A2(n391), .B0(n173), .Y(n383) );
  BUFX2 U684 ( .A(n358), .Y(n124) );
  NAND4X1 U685 ( .A(n771), .B(n597), .C(n772), .D(n762), .Y(n768) );
  NAND4X1 U686 ( .A(n1090), .B(n948), .C(n1091), .D(n1081), .Y(n1087) );
  NAND4X1 U687 ( .A(n669), .B(n788), .C(n581), .D(n837), .Y(n827) );
  AOI32X1 U688 ( .A0(n752), .A1(n77), .A2(n1637), .B0(n787), .B1(n75), .Y(n837) );
  NAND4X1 U689 ( .A(n1020), .B(n1107), .C(n932), .D(n1186), .Y(n1176) );
  AOI32X1 U690 ( .A0(n1071), .A1(n34), .A2(n1542), .B0(n1106), .B1(n36), .Y(
        n1186) );
  OAI31XL U691 ( .A0(n1614), .A1(n387), .A2(n388), .B0(n1596), .Y(n384) );
  NOR2X1 U692 ( .A(n361), .B(n348), .Y(n466) );
  OAI31XL U693 ( .A0(n398), .A1(n58), .A2(n196), .B0(n551), .Y(n550) );
  BUFX2 U694 ( .A(n1018), .Y(n146) );
  AOI2BB2X1 U695 ( .B0(n253), .B1(n1663), .A0N(n177), .A1N(n159), .Y(n833) );
  AOI2BB2X1 U696 ( .B0(n214), .B1(n1522), .A0N(n166), .A1N(n148), .Y(n1182) );
  BUFX2 U697 ( .A(n585), .Y(n155) );
  NOR2X1 U698 ( .A(n4), .B(n1582), .Y(n278) );
  OAI31XL U699 ( .A0(n747), .A1(n75), .A2(n87), .B0(n748), .Y(n746) );
  OAI21XL U700 ( .A0(n744), .A1(n613), .B0(n1661), .Y(n748) );
  OAI31XL U701 ( .A0(n1066), .A1(n36), .A2(n28), .B0(n1067), .Y(n1065) );
  OAI21XL U702 ( .A0(n1063), .A1(n964), .B0(n1505), .Y(n1067) );
  NAND2X1 U703 ( .A(n115), .B(n1668), .Y(n587) );
  INVX1 U704 ( .A(n7), .Y(n46) );
  NAND2X1 U705 ( .A(n1664), .B(n223), .Y(n771) );
  NAND2X1 U706 ( .A(n1531), .B(n213), .Y(n1090) );
  NAND3BX1 U707 ( .AN(n399), .B(n400), .C(n401), .Y(n392) );
  OAI222XL U708 ( .A0(n402), .A1(n65), .B0(n361), .B1(n69), .C0(n403), .C1(
        n348), .Y(n399) );
  AOI2BB2X1 U709 ( .B0(n70), .B1(n79), .A0N(n253), .A1N(n160), .Y(n908) );
  AOI2BB2X1 U710 ( .B0(n37), .B1(n30), .A0N(n214), .A1N(n149), .Y(n1257) );
  BUFX2 U711 ( .A(n574), .Y(n158) );
  BUFX2 U712 ( .A(n925), .Y(n147) );
  NAND3BX1 U713 ( .AN(n1307), .B(n1308), .C(n1309), .Y(n1302) );
  AOI222XL U714 ( .A0(n49), .A1(n1574), .B0(n1581), .B1(n191), .C0(n1558), 
        .C1(n334), .Y(n1309) );
  NAND3BX1 U715 ( .AN(n625), .B(n626), .C(n627), .Y(n618) );
  OAI222XL U716 ( .A0(n628), .A1(n74), .B0(n587), .B1(n73), .C0(n629), .C1(
        n158), .Y(n625) );
  INVX1 U717 ( .A(n275), .Y(n1553) );
  OR4X1 U718 ( .A(n724), .B(n744), .C(n616), .D(n730), .Y(n741) );
  OR4X1 U719 ( .A(n1043), .B(n1063), .C(n967), .D(n1049), .Y(n1060) );
  INVX1 U720 ( .A(n354), .Y(n1603) );
  AO21X1 U721 ( .A0(n249), .A1(n284), .B0(n51), .Y(n268) );
  NAND4BX1 U722 ( .AN(n852), .B(n598), .C(n594), .D(n853), .Y(n849) );
  AOI222XL U723 ( .A0(n76), .A1(n187), .B0(n253), .B1(n854), .C0(n773), .C1(
        n75), .Y(n853) );
  NAND2X1 U724 ( .A(n721), .B(n668), .Y(n854) );
  NAND4BX1 U725 ( .AN(n1201), .B(n949), .C(n945), .D(n1202), .Y(n1198) );
  AOI222XL U726 ( .A0(n33), .A1(n184), .B0(n214), .B1(n1203), .C0(n1092), .C1(
        n36), .Y(n1202) );
  NAND2X1 U727 ( .A(n1040), .B(n1019), .Y(n1203) );
  OAI221XL U728 ( .A0(n186), .A1(n575), .B0(sboxw[25]), .B1(n162), .C0(n833), 
        .Y(n831) );
  OAI221XL U729 ( .A0(n182), .A1(n152), .B0(sboxw[17]), .B1(n151), .C0(n1182), 
        .Y(n1180) );
  BUFX2 U730 ( .A(n645), .Y(n156) );
  BUFX2 U731 ( .A(n622), .Y(n162) );
  BUFX2 U732 ( .A(n973), .Y(n151) );
  BUFX2 U733 ( .A(n996), .Y(n145) );
  BUFX2 U734 ( .A(n951), .Y(n150) );
  BUFX2 U735 ( .A(n936), .Y(n144) );
  OAI31XL U736 ( .A0(n275), .A1(n49), .A2(n45), .B0(n1377), .Y(n1376) );
  OAI21XL U737 ( .A0(n338), .A1(n330), .B0(n6), .Y(n1377) );
  NAND4BX1 U738 ( .AN(n604), .B(n598), .C(n588), .D(n723), .Y(n718) );
  AOI211X1 U739 ( .A0(n1656), .A1(n1642), .B0(n724), .C0(n725), .Y(n723) );
  AOI2BB1X1 U740 ( .A0N(n1662), .A1N(n76), .B0(n157), .Y(n725) );
  NAND4BX1 U741 ( .AN(n955), .B(n949), .C(n939), .D(n1042), .Y(n1037) );
  AOI211X1 U742 ( .A0(n1513), .A1(n40), .B0(n1043), .C0(n1044), .Y(n1042) );
  AOI2BB1X1 U743 ( .A0N(n1514), .A1N(n33), .B0(n1018), .Y(n1044) );
  BUFX2 U744 ( .A(n594), .Y(n160) );
  BUFX2 U745 ( .A(n945), .Y(n149) );
  OAI22XL U746 ( .A0(n797), .A1(n635), .B0(n798), .B1(n633), .Y(n796) );
  AOI211X1 U747 ( .A0(n1645), .A1(n81), .B0(n800), .C0(n801), .Y(n797) );
  AOI221XL U748 ( .A0(n1663), .A1(n219), .B0(n71), .B1(n1664), .C0(n799), .Y(
        n798) );
  OAI22XL U749 ( .A0(n622), .A1(n155), .B0(n218), .B1(n159), .Y(n801) );
  INVX1 U750 ( .A(n407), .Y(n1590) );
  BUFX2 U751 ( .A(n1072), .Y(n148) );
  AOI211X1 U752 ( .A0(n1504), .A1(n182), .B0(n1245), .C0(n1246), .Y(n1236) );
  OAI31XL U753 ( .A0(n975), .A1(n1517), .A2(n182), .B0(n1190), .Y(n1246) );
  OAI222XL U754 ( .A0(n35), .A1(n958), .B0(n37), .B1(n1193), .C0(n1247), .C1(
        n165), .Y(n1245) );
  NOR4X1 U755 ( .A(n1248), .B(n1249), .C(n1528), .D(n1201), .Y(n1247) );
  AOI211X1 U756 ( .A0(n326), .A1(n1586), .B0(n1449), .C0(n1578), .Y(n1448) );
  INVX1 U757 ( .A(n674), .Y(n1645) );
  INVX1 U758 ( .A(n1025), .Y(n1538) );
  OAI2BB1X1 U759 ( .A0N(n1596), .A1N(n473), .B0(n381), .Y(n471) );
  INVX1 U760 ( .A(n747), .Y(n1659) );
  NAND2X1 U761 ( .A(n910), .B(n574), .Y(n895) );
  XOR2X1 U762 ( .A(n77), .B(n218), .Y(n910) );
  NAND2X1 U763 ( .A(n1259), .B(n925), .Y(n1244) );
  XOR2X1 U764 ( .A(n34), .B(n208), .Y(n1259) );
  INVX1 U765 ( .A(n682), .Y(n1644) );
  INVX1 U766 ( .A(n1033), .Y(n1539) );
  INVX1 U767 ( .A(n624), .Y(n1666) );
  OAI221XL U768 ( .A0(n48), .A1(n258), .B0(n52), .B1(n138), .C0(n1567), .Y(
        n324) );
  INVX1 U769 ( .A(n328), .Y(n1567) );
  AO22X1 U770 ( .A0(n1597), .A1(n1615), .B0(n1596), .B1(n388), .Y(n394) );
  OAI222XL U771 ( .A0(n66), .A1(n131), .B0(n124), .B1(n495), .C0(n494), .C1(
        n456), .Y(n556) );
  INVX1 U772 ( .A(n119), .Y(n86) );
  INVX1 U773 ( .A(sboxw[20]), .Y(n27) );
  OAI222XL U774 ( .A0(sboxw[25]), .A1(n668), .B0(n157), .B1(n587), .C0(n115), 
        .C1(n840), .Y(n882) );
  OAI222XL U775 ( .A0(sboxw[17]), .A1(n1019), .B0(n146), .B1(n938), .C0(n107), 
        .C1(n1189), .Y(n1231) );
  OAI2BB1X1 U776 ( .A0N(n6), .A1N(n1369), .B0(n297), .Y(n1362) );
  OAI21XL U777 ( .A0(n48), .A1(n1582), .B0(n191), .Y(n1369) );
  OAI222XL U778 ( .A0(n48), .A1(n297), .B0(n171), .B1(n311), .C0(n312), .C1(
        n169), .Y(n308) );
  NOR4X1 U779 ( .A(n313), .B(n314), .C(n1572), .D(n315), .Y(n312) );
  OAI21XL U780 ( .A0(n189), .A1(n316), .B0(n317), .Y(n314) );
  OAI222XL U781 ( .A0(n49), .A1(n138), .B0(n139), .B1(n10), .C0(n172), .C1(
        n133), .Y(n313) );
  OAI222XL U782 ( .A0(n74), .A1(n607), .B0(n71), .B1(n844), .C0(n898), .C1(
        n180), .Y(n896) );
  NOR4X1 U783 ( .A(n899), .B(n900), .C(n1635), .D(n852), .Y(n898) );
  OAI222XL U784 ( .A0(n75), .A1(n159), .B0(n73), .B1(n575), .C0(n1637), .C1(
        n622), .Y(n899) );
  OAI21XL U785 ( .A0(n585), .A1(n629), .B0(n679), .Y(n900) );
  AO22X1 U786 ( .A0(n168), .A1(n1569), .B0(n6), .B1(n1298), .Y(n1304) );
  OAI222XL U787 ( .A0(n139), .A1(n192), .B0(n136), .B1(n305), .C0(n288), .C1(
        n51), .Y(n300) );
  BUFX2 U788 ( .A(n4), .Y(n191) );
  AOI222XL U789 ( .A0(n65), .A1(n1624), .B0(n515), .B1(n196), .C0(n1609), .C1(
        n128), .Y(n545) );
  AOI211X1 U790 ( .A0(n664), .A1(n87), .B0(n665), .C0(n666), .Y(n662) );
  OAI22XL U791 ( .A0(n161), .A1(n667), .B0(n223), .B1(n594), .Y(n666) );
  OAI221XL U792 ( .A0(n584), .A1(n668), .B0(n219), .B1(n649), .C0(n669), .Y(
        n665) );
  AOI211X1 U793 ( .A0(n69), .A1(n60), .B0(n694), .C0(n695), .Y(n689) );
  OAI22XL U794 ( .A0(n21), .A1(n129), .B0(n15), .B1(n402), .Y(n695) );
  OAI221XL U795 ( .A0(n1610), .A1(n128), .B0(n199), .B1(n403), .C0(n696), .Y(
        n694) );
  AOI211X1 U796 ( .A0(n1015), .A1(n28), .B0(n1016), .C0(n1017), .Y(n1013) );
  OAI22XL U797 ( .A0(n951), .A1(n146), .B0(n213), .B1(n149), .Y(n1017) );
  OAI221XL U798 ( .A0(n142), .A1(n1019), .B0(n209), .B1(n1000), .C0(n1020), 
        .Y(n1016) );
  BUFX2 U799 ( .A(n753), .Y(n159) );
  BUFX2 U800 ( .A(n4), .Y(n192) );
  INVX1 U801 ( .A(n119), .Y(n87) );
  AOI221XL U802 ( .A0(n1592), .A1(n536), .B0(n1591), .B1(n537), .C0(n538), .Y(
        n535) );
  NAND4BX1 U803 ( .AN(n389), .B(n530), .C(n546), .D(n547), .Y(n536) );
  OAI22XL U804 ( .A0(n539), .A1(n409), .B0(n540), .B1(n407), .Y(n538) );
  OAI31XL U805 ( .A0(n4), .A1(n46), .A2(n47), .B0(n1287), .Y(n1286) );
  OAI31XL U806 ( .A0(n295), .A1(n50), .A2(n1563), .B0(n310), .Y(n309) );
  OAI31XL U807 ( .A0(n58), .A1(n69), .A2(n353), .B0(n445), .Y(n707) );
  OAI31XL U808 ( .A0(n624), .A1(n1667), .A2(n186), .B0(n841), .Y(n897) );
  INVX1 U809 ( .A(n273), .Y(n1576) );
  AOI211X1 U810 ( .A0(n378), .A1(n1600), .B0(n379), .C0(n380), .Y(n341) );
  OAI22XL U811 ( .A0(n24), .A1(n381), .B0(n382), .B1(n1597), .Y(n380) );
  NAND4X1 U812 ( .A(n383), .B(n384), .C(n385), .D(n386), .Y(n379) );
  AOI211X1 U813 ( .A0(n1607), .A1(n124), .B0(n11), .C0(n1617), .Y(n382) );
  OAI211X1 U814 ( .A0(n1644), .A1(n645), .B0(n1665), .C0(n678), .Y(n658) );
  INVX1 U815 ( .A(n681), .Y(n1665) );
  NOR2BX1 U816 ( .AN(n679), .B(n680), .Y(n678) );
  OAI211X1 U817 ( .A0(n1539), .A1(n996), .B0(n1532), .C0(n1029), .Y(n1009) );
  INVX1 U818 ( .A(n1032), .Y(n1532) );
  NOR2BX1 U819 ( .AN(n1030), .B(n1031), .Y(n1029) );
  OAI211X1 U820 ( .A0(sboxw[25]), .A1(n657), .B0(n669), .C0(n833), .Y(n848) );
  OAI211X1 U821 ( .A0(sboxw[17]), .A1(n1008), .B0(n1020), .C0(n1182), .Y(n1197) );
  OAI211X1 U822 ( .A0(n71), .A1(n657), .B0(n772), .C0(n783), .Y(n782) );
  OAI211X1 U823 ( .A0(n38), .A1(n1008), .B0(n1091), .C0(n1102), .Y(n1101) );
  OAI211X1 U824 ( .A0(n188), .A1(n629), .B0(n679), .C0(n802), .Y(n800) );
  AOI2BB2X1 U825 ( .B0(n1652), .B1(n218), .A0N(n584), .A1N(n628), .Y(n802) );
  OAI211X1 U826 ( .A0(n184), .A1(n980), .B0(n1030), .C0(n1151), .Y(n1149) );
  AOI2BB2X1 U827 ( .B0(n1518), .B1(n208), .A0N(n142), .A1N(n979), .Y(n1151) );
  OAI22XL U828 ( .A0(n131), .A1(n16), .B0(n193), .B1(n495), .Y(n543) );
  OAI211X1 U829 ( .A0(n15), .A1(n403), .B0(n453), .C0(n544), .Y(n542) );
  INVX1 U830 ( .A(n770), .Y(n1650) );
  INVX1 U831 ( .A(n1089), .Y(n1536) );
  INVX1 U832 ( .A(n1287), .Y(n1557) );
  INVX1 U833 ( .A(n840), .Y(n1641) );
  INVX1 U834 ( .A(n1189), .Y(n1537) );
  INVX1 U835 ( .A(n305), .Y(n1555) );
  OAI22XL U836 ( .A0(n586), .A1(n721), .B0(n784), .B1(n602), .Y(n864) );
  OAI22XL U837 ( .A0(n937), .A1(n1040), .B0(n1103), .B1(n953), .Y(n1213) );
  OAI22XL U838 ( .A0(n71), .A1(n851), .B0(n865), .B1(n1675), .Y(n862) );
  AOI2BB2X1 U839 ( .B0(n79), .B1(n219), .A0N(n622), .A1N(n73), .Y(n865) );
  OAI22XL U840 ( .A0(n38), .A1(n1200), .B0(n1214), .B1(n1506), .Y(n1211) );
  AOI2BB2X1 U841 ( .B0(n30), .B1(n209), .A0N(n973), .A1N(n39), .Y(n1214) );
  OAI2BB2XL U842 ( .B0(n157), .B1(n810), .A0N(n667), .A1N(n637), .Y(n863) );
  OAI2BB2XL U843 ( .B0(n1018), .B1(n1159), .A0N(n146), .A1N(n988), .Y(n1212)
         );
  NOR3X1 U844 ( .A(n747), .B(n72), .C(n721), .Y(n589) );
  NOR3X1 U845 ( .A(n1066), .B(n40), .C(n1040), .Y(n940) );
  OAI22XL U846 ( .A0(n150), .A1(n925), .B0(n144), .B1(n1019), .Y(n1093) );
  NOR2X1 U847 ( .A(n602), .B(n752), .Y(n818) );
  NOR2X1 U848 ( .A(n953), .B(n1071), .Y(n1167) );
  NAND2X1 U849 ( .A(n179), .B(n84), .Y(n635) );
  NAND2X1 U850 ( .A(n164), .B(n25), .Y(n986) );
  NAND2X1 U851 ( .A(n1662), .B(n223), .Y(n581) );
  NAND2X1 U852 ( .A(n1514), .B(n213), .Y(n932) );
  NAND2X1 U853 ( .A(n1531), .B(n208), .Y(n1020) );
  NAND4BX1 U854 ( .AN(n1347), .B(n285), .C(n1348), .D(n317), .Y(n1330) );
  NOR2X1 U855 ( .A(n600), .B(n747), .Y(n637) );
  NOR2X1 U856 ( .A(n150), .B(n1066), .Y(n988) );
  NAND2X1 U857 ( .A(n107), .B(n1534), .Y(n938) );
  NOR2X1 U858 ( .A(n156), .B(n223), .Y(n614) );
  NOR2X1 U859 ( .A(n145), .B(n213), .Y(n965) );
  NAND2X1 U860 ( .A(n223), .B(n637), .Y(n612) );
  NAND2X1 U861 ( .A(n213), .B(n988), .Y(n963) );
  NAND3BX1 U862 ( .AN(n976), .B(n977), .C(n978), .Y(n969) );
  OAI222XL U863 ( .A0(n979), .A1(n35), .B0(n938), .B1(n39), .C0(n980), .C1(
        n147), .Y(n976) );
  BUFX2 U864 ( .A(n667), .Y(n157) );
  BUFX2 U865 ( .A(n600), .Y(n161) );
  INVX1 U866 ( .A(n1066), .Y(n1509) );
  NAND2X1 U867 ( .A(n787), .B(n218), .Y(n836) );
  NAND2X1 U868 ( .A(n1106), .B(n208), .Y(n1185) );
  OAI2BB1X1 U869 ( .A0N(n424), .A1N(n19), .B0(n124), .Y(n527) );
  INVX1 U870 ( .A(n975), .Y(n1502) );
  NAND2X1 U871 ( .A(n818), .B(n223), .Y(n841) );
  NAND2X1 U872 ( .A(n1167), .B(n213), .Y(n1190) );
  BUFX2 U873 ( .A(n1675), .Y(n180) );
  INVX1 U874 ( .A(sboxw[20]), .Y(n28) );
  INVX1 U875 ( .A(n1313), .Y(n1545) );
  INVX1 U876 ( .A(n633), .Y(n1672) );
  INVX1 U877 ( .A(n984), .Y(n1345) );
  OAI21XL U878 ( .A0(n1414), .A1(n1415), .B0(n1543), .Y(n1413) );
  OAI31XL U879 ( .A0(n1427), .A1(n1428), .A2(n1429), .B0(n1544), .Y(n1412) );
  NOR4BBX1 U880 ( .AN(n1430), .BN(n1306), .C(n1436), .D(n1437), .Y(n1411) );
  NAND2X1 U881 ( .A(n100), .B(n169), .Y(n295) );
  OAI22XL U882 ( .A0(n98), .A1(n100), .B0(n99), .B1(n140), .Y(n1321) );
  OAI22XL U883 ( .A0(n47), .A1(n206), .B0(n100), .B1(n140), .Y(n1342) );
  OAI21XL U884 ( .A0(n1421), .A1(n1313), .B0(n1422), .Y(n1414) );
  OAI31XL U885 ( .A0(n1423), .A1(n1424), .A2(n1425), .B0(n1546), .Y(n1422) );
  NAND2X1 U886 ( .A(n102), .B(n47), .Y(n258) );
  NAND2X1 U887 ( .A(sboxw[12]), .B(sboxw[10]), .Y(n281) );
  NAND2X1 U888 ( .A(n103), .B(n1582), .Y(n7) );
  NOR2X1 U889 ( .A(n99), .B(n102), .Y(n323) );
  NAND2X1 U890 ( .A(n1549), .B(sboxw[11]), .Y(n239) );
  NOR3X1 U891 ( .A(n236), .B(n1563), .C(n205), .Y(n1428) );
  NAND2X1 U892 ( .A(n9), .B(n100), .Y(n244) );
  AND2X2 U893 ( .A(sboxw[12]), .B(n1582), .Y(n9) );
  NAND2X1 U894 ( .A(n103), .B(n102), .Y(n287) );
  NAND2X1 U895 ( .A(n102), .B(n1568), .Y(n261) );
  OAI211X1 U896 ( .A0(n206), .A1(n239), .B0(n1368), .C0(n1438), .Y(n1436) );
  INVX1 U897 ( .A(n102), .Y(n1582) );
  INVX1 U898 ( .A(sboxw[10]), .Y(n47) );
  BUFX2 U899 ( .A(n334), .Y(n140) );
  INVX1 U900 ( .A(sboxw[14]), .Y(n41) );
  OAI22XL U901 ( .A0(n90), .A1(n193), .B0(n64), .B1(n348), .Y(n456) );
  OAI21XL U902 ( .A0(n198), .A1(n19), .B0(n131), .Y(n455) );
  NAND2X1 U903 ( .A(n68), .B(n91), .Y(n700) );
  OAI22XL U904 ( .A0(n54), .A1(n435), .B0(n436), .B1(n437), .Y(n434) );
  AOI211X1 U905 ( .A0(n438), .A1(n58), .B0(n439), .C0(n440), .Y(n436) );
  OAI22XL U906 ( .A0(n19), .A1(n441), .B0(n198), .B1(n368), .Y(n440) );
  OAI221XL U907 ( .A0(n123), .A1(n442), .B0(n194), .B1(n423), .C0(n443), .Y(
        n439) );
  AOI2BB2X1 U908 ( .B0(n63), .B1(n18), .A0N(n200), .A1N(n63), .Y(n22) );
  NAND2X1 U909 ( .A(n106), .B(n41), .Y(n1313) );
  NAND4X1 U910 ( .A(n447), .B(n445), .C(n446), .D(n444), .Y(n433) );
  OAI21XL U911 ( .A0(n1614), .A1(n1626), .B0(n1600), .Y(n446) );
  AOI222XL U912 ( .A0(n56), .A1(n448), .B0(n94), .B1(n449), .C0(n450), .C1(
        n173), .Y(n447) );
  NAND2X1 U913 ( .A(n90), .B(n61), .Y(n431) );
  NAND2X1 U914 ( .A(sboxw[4]), .B(n91), .Y(n17) );
  NAND2X1 U915 ( .A(n193), .B(n198), .Y(n358) );
  INVX1 U916 ( .A(n18), .Y(n348) );
  AOI2BB2X1 U917 ( .B0(n67), .B1(n1619), .A0N(n199), .A1N(n368), .Y(n1491) );
  NAND2X1 U918 ( .A(n1621), .B(n198), .Y(n513) );
  INVX1 U919 ( .A(sboxw[3]), .Y(n1623) );
  INVX1 U920 ( .A(n92), .Y(n57) );
  NAND2X1 U921 ( .A(n92), .B(n1623), .Y(n494) );
  BUFX2 U922 ( .A(n197), .Y(n195) );
  NAND2X1 U923 ( .A(n91), .B(n57), .Y(n419) );
  NAND2X1 U924 ( .A(n55), .B(n89), .Y(n368) );
  NAND2X1 U925 ( .A(n90), .B(n8), .Y(n396) );
  AND2X2 U926 ( .A(n92), .B(n91), .Y(n8) );
  NAND2X1 U927 ( .A(n89), .B(n1607), .Y(n495) );
  NAND2X1 U928 ( .A(n198), .B(n195), .Y(n441) );
  NAND2X1 U929 ( .A(n200), .B(n195), .Y(n359) );
  AO21X1 U930 ( .A0(n201), .A1(n1605), .B0(n391), .Y(n449) );
  AOI221XL U931 ( .A0(n1598), .A1(n68), .B0(n66), .B1(n411), .C0(n412), .Y(
        n410) );
  OAI22XL U932 ( .A0(n93), .A1(n413), .B0(n414), .B1(n173), .Y(n412) );
  AOI211X1 U933 ( .A0(n1616), .A1(n20), .B0(n416), .C0(n417), .Y(n413) );
  INVX1 U934 ( .A(n93), .Y(n1597) );
  INVX1 U935 ( .A(n1350), .Y(n1544) );
  AOI211X1 U936 ( .A0(sboxw[13]), .A1(n1302), .B0(n1303), .C0(n1304), .Y(n1265) );
  NAND2X1 U937 ( .A(n93), .B(n53), .Y(n407) );
  NAND2X1 U938 ( .A(n1604), .B(n198), .Y(n354) );
  OAI222XL U939 ( .A0(sboxw[1]), .A1(n381), .B0(n94), .B1(n1474), .C0(n1475), 
        .C1(n173), .Y(n1472) );
  AOI211X1 U940 ( .A0(n1607), .A1(n1478), .B0(n390), .C0(n378), .Y(n1474) );
  OAI21XL U941 ( .A0(n1608), .A1(n430), .B0(n696), .Y(n1477) );
  NAND2X1 U942 ( .A(n1605), .B(n198), .Y(n355) );
  OAI22XL U943 ( .A0(n200), .A1(n423), .B0(n1630), .B1(n424), .Y(n422) );
  NOR3X1 U944 ( .A(n66), .B(n89), .C(n1608), .Y(n712) );
  NAND2X1 U945 ( .A(n94), .B(n64), .Y(n489) );
  NOR2X1 U946 ( .A(n64), .B(n91), .Y(n529) );
  NAND2X1 U947 ( .A(n89), .B(n92), .Y(n442) );
  NOR2X1 U948 ( .A(n431), .B(n200), .Y(n390) );
  AOI221XL U949 ( .A0(n1364), .A1(n168), .B0(n106), .B1(n1365), .C0(n1366), 
        .Y(n1363) );
  OAI21XL U950 ( .A0(n172), .A1(n316), .B0(n1367), .Y(n1366) );
  NAND2X1 U951 ( .A(n90), .B(n174), .Y(n398) );
  NAND2X1 U952 ( .A(n90), .B(n91), .Y(n424) );
  INVX1 U953 ( .A(n200), .Y(n199) );
  INVX1 U954 ( .A(n92), .Y(n58) );
  BUFX2 U955 ( .A(n197), .Y(n196) );
  INVX1 U956 ( .A(sboxw[6]), .Y(n54) );
  AOI222XL U957 ( .A0(n62), .A1(n199), .B0(n1598), .B1(n16), .C0(n93), .C1(
        n367), .Y(n366) );
  OAI211X1 U958 ( .A0(n201), .A1(n130), .B0(n369), .C0(n370), .Y(n367) );
  AND2X2 U959 ( .A(n371), .B(n372), .Y(n370) );
  NAND2X1 U960 ( .A(n1269), .B(n1543), .Y(n1268) );
  OAI211X1 U961 ( .A0(n1270), .A1(n229), .B0(n1271), .C0(n1272), .Y(n1269) );
  NOR4X1 U962 ( .A(n1290), .B(n1291), .C(n1564), .D(n1292), .Y(n1270) );
  OAI31XL U963 ( .A0(n1284), .A1(n1285), .A2(n1286), .B0(n1547), .Y(n1271) );
  OAI31XL U964 ( .A0(n1280), .A1(n1577), .A2(n1559), .B0(sboxw[13]), .Y(n1279)
         );
  INVX1 U965 ( .A(n1282), .Y(n1577) );
  OAI31XL U966 ( .A0(n1273), .A1(n1274), .A2(n1275), .B0(n42), .Y(n1272) );
  OAI22XL U967 ( .A0(n287), .A1(n1276), .B0(n189), .B1(n1277), .Y(n1275) );
  OAI221XL U968 ( .A0(n1586), .A1(n269), .B0(n206), .B1(n252), .C0(n1279), .Y(
        n1273) );
  AOI31X1 U969 ( .A0(n1629), .A1(sboxw[2]), .A2(n1608), .B0(n351), .Y(n350) );
  OAI31XL U970 ( .A0(n21), .A1(n353), .A2(n58), .B0(n354), .Y(n351) );
  INVX1 U971 ( .A(n95), .Y(n53) );
  INVX1 U972 ( .A(n1113), .Y(n1591) );
  AOI211X1 U973 ( .A0(n54), .A1(n1126), .B0(n1127), .C0(n1128), .Y(n1110) );
  OAI22XL U974 ( .A0(n170), .A1(n241), .B0(n242), .B1(n168), .Y(n232) );
  AOI221XL U975 ( .A0(n240), .A1(n1586), .B0(n1551), .B1(n190), .C0(n1317), 
        .Y(n1316) );
  AOI221XL U976 ( .A0(n1570), .A1(n140), .B0(n1574), .B1(n205), .C0(n1325), 
        .Y(n1314) );
  AOI2BB2X1 U977 ( .B0(n67), .B1(n1596), .A0N(n66), .A1N(n398), .Y(n395) );
  OAI222XL U978 ( .A0(n507), .A1(n173), .B0(n508), .B1(n489), .C0(n509), .C1(
        n93), .Y(n498) );
  AOI211X1 U979 ( .A0(n515), .A1(n194), .B0(n516), .C0(n1621), .Y(n507) );
  AOI222XL U980 ( .A0(n522), .A1(n93), .B0(n1596), .B1(n523), .C0(n524), .C1(
        n1597), .Y(n519) );
  NAND4X1 U981 ( .A(n528), .B(n427), .C(n527), .D(n442), .Y(n522) );
  AOI222XL U982 ( .A0(sboxw[13]), .A1(n1403), .B0(n6), .B1(n1404), .C0(n1405), 
        .C1(n168), .Y(n1400) );
  OAI221XL U983 ( .A0(n171), .A1(n244), .B0(n136), .B1(n133), .C0(n246), .Y(
        n1405) );
  NAND4X1 U984 ( .A(n1341), .B(n1339), .C(n1340), .D(n1338), .Y(n1331) );
  OAI21XL U985 ( .A0(n1283), .A1(n278), .B0(n1553), .Y(n1340) );
  NAND2X1 U986 ( .A(n1549), .B(n1346), .Y(n1338) );
  AOI222XL U987 ( .A0(n44), .A1(n1342), .B0(n105), .B1(n1343), .C0(n1344), 
        .C1(n168), .Y(n1341) );
  OAI222XL U988 ( .A0(sboxw[1]), .A1(n442), .B0(n441), .B1(n361), .C0(n63), 
        .C1(n700), .Y(n1137) );
  AOI2BB2X1 U989 ( .B0(n6), .B1(n170), .A0N(n170), .A1N(n295), .Y(n1305) );
  OAI222XL U990 ( .A0(n274), .A1(n275), .B0(n276), .B1(n168), .C0(n277), .C1(
        n106), .Y(n262) );
  AOI221XL U991 ( .A0(n46), .A1(n52), .B0(n1562), .B1(n135), .C0(n286), .Y(
        n274) );
  OAI222XL U992 ( .A0(n1392), .A1(n169), .B0(n1393), .B1(n275), .C0(sboxw[13]), 
        .C1(n1394), .Y(n1383) );
  OAI22XL U993 ( .A0(n42), .A1(n296), .B0(n1333), .B1(n229), .Y(n1332) );
  OAI221XL U994 ( .A0(n191), .A1(n281), .B0(sboxw[8]), .B1(n249), .C0(n1336), 
        .Y(n1335) );
  NAND2X1 U995 ( .A(n105), .B(n47), .Y(n275) );
  OAI31XL U996 ( .A0(n389), .A1(n1618), .A2(n472), .B0(n94), .Y(n1135) );
  AOI221XL U997 ( .A0(n1613), .A1(n194), .B0(n67), .B1(n1621), .C0(n541), .Y(
        n540) );
  NOR3X1 U998 ( .A(n170), .B(n100), .C(n1563), .Y(n315) );
  OAI22XL U999 ( .A0(n829), .A1(n663), .B0(n830), .B1(n635), .Y(n828) );
  AOI211X1 U1000 ( .A0(n73), .A1(n80), .B0(n834), .C0(n835), .Y(n829) );
  NOR4BX1 U1001 ( .AN(n788), .B(n831), .C(n832), .D(n1635), .Y(n830) );
  OAI221XL U1002 ( .A0(n1653), .A1(n574), .B0(n253), .B1(n629), .C0(n836), .Y(
        n834) );
  OAI22XL U1003 ( .A0(n1178), .A1(n1014), .B0(n1179), .B1(n986), .Y(n1177) );
  AOI211X1 U1004 ( .A0(n39), .A1(n31), .B0(n1183), .C0(n1184), .Y(n1178) );
  NOR4BX1 U1005 ( .AN(n1107), .B(n1180), .C(n1181), .D(n1528), .Y(n1179) );
  OAI221XL U1006 ( .A0(n1519), .A1(n925), .B0(n214), .B1(n980), .C0(n1185), 
        .Y(n1183) );
  AOI222XL U1007 ( .A0(n62), .A1(n175), .B0(n194), .B1(n1131), .C0(n1123), 
        .C1(n23), .Y(n1130) );
  AOI222XL U1008 ( .A0(n69), .A1(n1607), .B0(n1605), .B1(n196), .C0(n59), .C1(
        n359), .Y(n1129) );
  OAI22XL U1009 ( .A0(n106), .A1(n1318), .B0(n1319), .B1(n104), .Y(n1317) );
  OAI221XL U1010 ( .A0(n259), .A1(n140), .B0(n249), .B1(n141), .C0(n1324), .Y(
        n1322) );
  NAND2X1 U1011 ( .A(n1664), .B(n221), .Y(n598) );
  NAND2X1 U1012 ( .A(n1531), .B(n211), .Y(n949) );
  OAI211X1 U1013 ( .A0(n130), .A1(n123), .B0(n1606), .C0(n501), .Y(n500) );
  AOI221XL U1014 ( .A0(n1604), .A1(n18), .B0(n1616), .B1(n1630), .C0(n502), 
        .Y(n501) );
  NOR3X1 U1015 ( .A(n482), .B(n89), .C(n23), .Y(n502) );
  AOI2BB2X1 U1016 ( .B0(n200), .B1(n59), .A0N(n24), .A1N(n495), .Y(n400) );
  NAND3X1 U1017 ( .A(n90), .B(n441), .C(n1608), .Y(n505) );
  AOI222XL U1018 ( .A0(n1605), .A1(n359), .B0(n1625), .B1(n199), .C0(n1609), 
        .C1(n1630), .Y(n506) );
  NAND2X1 U1019 ( .A(n1599), .B(n200), .Y(n385) );
  NOR3X1 U1020 ( .A(n70), .B(sboxw[26]), .C(n1667), .Y(n852) );
  NOR3X1 U1021 ( .A(n37), .B(n108), .C(n1517), .Y(n1201) );
  NOR2X1 U1022 ( .A(n77), .B(sboxw[27]), .Y(n787) );
  NOR2X1 U1023 ( .A(n34), .B(sboxw[19]), .Y(n1106) );
  NAND2X1 U1024 ( .A(n1579), .B(n203), .Y(n273) );
  AOI221XL U1025 ( .A0(n1573), .A1(n191), .B0(n190), .B1(n1580), .C0(n271), 
        .Y(n270) );
  AOI221XL U1026 ( .A0(n49), .A1(n240), .B0(n1546), .B1(n1398), .C0(n1399), 
        .Y(n1381) );
  OAI22XL U1027 ( .A0(n1400), .A1(n42), .B0(n1401), .B1(n1313), .Y(n1399) );
  NAND2X1 U1028 ( .A(n117), .B(n81), .Y(n657) );
  NAND2X1 U1029 ( .A(n109), .B(n32), .Y(n1008) );
  OAI22XL U1030 ( .A0(n161), .A1(n221), .B0(n70), .B1(n721), .Y(n884) );
  OAI22XL U1031 ( .A0(n777), .A1(n85), .B0(n778), .B1(n633), .Y(n776) );
  AOI221XL U1032 ( .A0(n1669), .A1(n186), .B0(n83), .B1(n154), .C0(n779), .Y(
        n778) );
  AOI222XL U1033 ( .A0(n120), .A1(n780), .B0(n1661), .B1(n781), .C0(n782), 
        .C1(n1675), .Y(n777) );
  OAI211X1 U1034 ( .A0(n352), .A1(n650), .B0(n588), .C0(n159), .Y(n779) );
  OAI22XL U1035 ( .A0(n1096), .A1(n1499), .B0(n1097), .B1(n984), .Y(n1095) );
  AOI221XL U1036 ( .A0(n1516), .A1(n182), .B0(n1523), .B1(n143), .C0(n1098), 
        .Y(n1097) );
  AOI222XL U1037 ( .A0(n112), .A1(n1099), .B0(n1505), .B1(n1100), .C0(n1101), 
        .C1(n165), .Y(n1096) );
  OAI211X1 U1038 ( .A0(n215), .A1(n1001), .B0(n939), .C0(n1072), .Y(n1098) );
  OAI22XL U1039 ( .A0(n1146), .A1(n986), .B0(n1147), .B1(n984), .Y(n1145) );
  AOI221XL U1040 ( .A0(n1522), .A1(n209), .B0(n38), .B1(n1531), .C0(n1148), 
        .Y(n1147) );
  AOI211X1 U1041 ( .A0(n1538), .A1(n32), .B0(n1149), .C0(n1150), .Y(n1146) );
  OAI31XL U1042 ( .A0(n1535), .A1(n111), .A2(n147), .B0(n1055), .Y(n1148) );
  OAI22XL U1043 ( .A0(n118), .A1(n75), .B0(n1645), .B1(n161), .Y(n676) );
  OAI22XL U1044 ( .A0(n110), .A1(n36), .B0(n1538), .B1(n150), .Y(n1027) );
  NOR4BX1 U1045 ( .AN(n772), .B(n866), .C(n867), .D(n1655), .Y(n859) );
  OAI22XL U1046 ( .A0(n220), .A1(n649), .B0(n71), .B1(n1653), .Y(n867) );
  OAI222XL U1047 ( .A0(n157), .A1(n159), .B0(n578), .B1(n629), .C0(n657), .C1(
        n585), .Y(n866) );
  NOR4BX1 U1048 ( .AN(n1091), .B(n1215), .C(n1216), .D(n1512), .Y(n1208) );
  OAI22XL U1049 ( .A0(n210), .A1(n1000), .B0(n38), .B1(n1519), .Y(n1216) );
  OAI222XL U1050 ( .A0(n1018), .A1(n1072), .B0(n183), .B1(n980), .C0(n1008), 
        .C1(n144), .Y(n1215) );
  NOR4X1 U1051 ( .A(n487), .B(n488), .C(n1603), .D(n363), .Y(n457) );
  OAI31XL U1052 ( .A0(n489), .A1(n18), .A2(n58), .B0(n490), .Y(n488) );
  OAI222XL U1053 ( .A0(n381), .A1(n124), .B0(n93), .B1(n491), .C0(n492), .C1(
        n173), .Y(n487) );
  OAI21XL U1054 ( .A0(n486), .A1(n387), .B0(n1596), .Y(n490) );
  NAND2X1 U1055 ( .A(n1593), .B(n91), .Y(n552) );
  AOI2BB2X1 U1056 ( .B0(n266), .B1(n79), .A0N(n187), .A1N(n159), .Y(n626) );
  AOI2BB2X1 U1057 ( .B0(n216), .B1(n30), .A0N(n184), .A1N(n148), .Y(n977) );
  AOI2BB2X1 U1058 ( .B0(n153), .B1(n117), .A0N(n116), .A1N(n74), .Y(n586) );
  AOI2BB2X1 U1059 ( .B0(n142), .B1(n109), .A0N(n108), .A1N(n35), .Y(n937) );
  NAND4X1 U1060 ( .A(n1388), .B(n1389), .C(n1390), .D(n1391), .Y(n1384) );
  AOI222XL U1061 ( .A0(n1560), .A1(n5), .B0(n1584), .B1(n204), .C0(n1564), 
        .C1(n1587), .Y(n1391) );
  AOI2BB2X1 U1062 ( .B0(n118), .B1(n253), .A0N(n253), .A1N(n752), .Y(n784) );
  AOI2BB2X1 U1063 ( .B0(n110), .B1(n214), .A0N(n214), .A1N(n1071), .Y(n1103)
         );
  NAND2X1 U1064 ( .A(sboxw[27]), .B(n115), .Y(n770) );
  NAND2X1 U1065 ( .A(sboxw[19]), .B(n107), .Y(n1089) );
  NAND2X1 U1066 ( .A(n116), .B(n179), .Y(n624) );
  OAI211X1 U1067 ( .A0(n21), .A1(n552), .B0(n553), .C0(n554), .Y(n548) );
  OAI21XL U1068 ( .A0(n387), .A1(n1621), .B0(n1597), .Y(n553) );
  OAI21XL U1069 ( .A0(n555), .A1(n556), .B0(n93), .Y(n554) );
  OAI222XL U1070 ( .A0(n607), .A1(n154), .B0(n120), .B1(n749), .C0(n750), .C1(
        n180), .Y(n745) );
  AOI211X1 U1071 ( .A0(n1642), .A1(n79), .B0(n751), .C0(n1634), .Y(n750) );
  OA21XL U1072 ( .A0(n752), .A1(n155), .B0(n626), .Y(n749) );
  OAI22XL U1073 ( .A0(n260), .A1(n645), .B0(n72), .B1(n622), .Y(n751) );
  OAI222XL U1074 ( .A0(n958), .A1(n143), .B0(n112), .B1(n1068), .C0(n1069), 
        .C1(n165), .Y(n1064) );
  AOI211X1 U1075 ( .A0(n40), .A1(n30), .B0(n1070), .C0(n1521), .Y(n1069) );
  OA21XL U1076 ( .A0(n1071), .A1(n936), .B0(n977), .Y(n1068) );
  OAI22XL U1077 ( .A0(n215), .A1(n996), .B0(n40), .B1(n973), .Y(n1070) );
  NOR4X1 U1078 ( .A(n869), .B(n870), .C(n617), .D(n1643), .Y(n857) );
  OAI32X1 U1079 ( .A0(n222), .A1(sboxw[28]), .A2(n116), .B0(n73), .B1(n770), 
        .Y(n870) );
  OAI222XL U1080 ( .A0(n657), .A1(n584), .B0(n155), .B1(n649), .C0(n186), .C1(
        n645), .Y(n869) );
  NOR4X1 U1081 ( .A(n1218), .B(n1219), .C(n968), .D(n1520), .Y(n1206) );
  OAI32X1 U1082 ( .A0(n212), .A1(n111), .A2(n108), .B0(n39), .B1(n1089), .Y(
        n1219) );
  OAI222XL U1083 ( .A0(n1008), .A1(n142), .B0(n936), .B1(n1000), .C0(n182), 
        .C1(n996), .Y(n1218) );
  AOI22X1 U1084 ( .A0(n734), .A1(n179), .B0(n121), .B1(n735), .Y(n733) );
  OAI21XL U1085 ( .A0(n218), .A1(n650), .B0(n162), .Y(n735) );
  OAI21XL U1086 ( .A0(n75), .A1(n645), .B0(n736), .Y(n734) );
  AOI22X1 U1087 ( .A0(n1053), .A1(n164), .B0(n113), .B1(n1054), .Y(n1052) );
  OAI21XL U1088 ( .A0(n208), .A1(n1001), .B0(n151), .Y(n1054) );
  OAI21XL U1089 ( .A0(n36), .A1(n145), .B0(n1055), .Y(n1053) );
  NAND2X1 U1090 ( .A(n323), .B(n98), .Y(n304) );
  OAI21XL U1091 ( .A0(n483), .A1(n484), .B0(n94), .Y(n480) );
  OR4X1 U1092 ( .A(n466), .B(n486), .C(n390), .D(n472), .Y(n483) );
  OAI21XL U1093 ( .A0(n1373), .A1(n1374), .B0(n106), .Y(n1371) );
  NAND4BBXL U1094 ( .AN(n307), .BN(n338), .C(n1357), .D(n302), .Y(n1373) );
  NAND2X1 U1095 ( .A(n72), .B(n118), .Y(n840) );
  NAND2X1 U1096 ( .A(n1541), .B(n110), .Y(n1189) );
  NAND2X1 U1097 ( .A(n203), .B(n1558), .Y(n1287) );
  OAI31XL U1098 ( .A0(n431), .A1(n93), .A2(n194), .B0(n377), .Y(n1116) );
  OAI31XL U1099 ( .A0(n244), .A1(sboxw[8]), .A2(sboxw[13]), .B0(n245), .Y(n231) );
  NAND4BX1 U1100 ( .AN(n589), .B(n590), .C(n591), .D(n592), .Y(n570) );
  AOI2BB2X1 U1101 ( .B0(n599), .B1(n154), .A0N(n161), .A1N(n601), .Y(n591) );
  NAND3X1 U1102 ( .A(n185), .B(n1668), .C(n1666), .Y(n590) );
  AOI222XL U1103 ( .A0(n76), .A1(n253), .B0(n1657), .B1(n585), .C0(n120), .C1(
        n593), .Y(n592) );
  NAND4BX1 U1104 ( .AN(n940), .B(n941), .C(n942), .D(n943), .Y(n921) );
  AOI2BB2X1 U1105 ( .B0(n950), .B1(n143), .A0N(n951), .A1N(n952), .Y(n942) );
  NAND3X1 U1106 ( .A(n181), .B(n1534), .C(n1502), .Y(n941) );
  AOI222XL U1107 ( .A0(n33), .A1(n214), .B0(n1507), .B1(n144), .C0(n112), .C1(
        n944), .Y(n943) );
  NAND4BX1 U1108 ( .AN(n680), .B(n761), .C(n161), .D(n803), .Y(n795) );
  AOI222XL U1109 ( .A0(n74), .A1(n1649), .B0(n773), .B1(n221), .C0(n1652), 
        .C1(n574), .Y(n803) );
  NAND4BX1 U1110 ( .AN(n1031), .B(n1080), .C(n951), .D(n1152), .Y(n1144) );
  AOI222XL U1111 ( .A0(n35), .A1(n1535), .B0(n1092), .B1(n210), .C0(n1518), 
        .C1(n925), .Y(n1152) );
  AOI2BB2X1 U1112 ( .B0(n123), .B1(sboxw[2]), .A0N(n90), .A1N(n65), .Y(n360)
         );
  AOI2BB2X1 U1113 ( .B0(n102), .B1(n204), .A0N(n204), .A1N(n7), .Y(n235) );
  NAND4X1 U1114 ( .A(n652), .B(n669), .C(n838), .D(n839), .Y(n826) );
  AOI22X1 U1115 ( .A0(n188), .A1(n787), .B0(n1641), .B1(n116), .Y(n838) );
  AOI222XL U1116 ( .A0(n83), .A1(n157), .B0(n1654), .B1(n260), .C0(n1656), 
        .C1(n154), .Y(n839) );
  NAND4X1 U1117 ( .A(n1003), .B(n1020), .C(n1187), .D(n1188), .Y(n1175) );
  AOI22X1 U1118 ( .A0(n184), .A1(n1106), .B0(n1537), .B1(n108), .Y(n1187) );
  AOI222XL U1119 ( .A0(n1523), .A1(n1018), .B0(n1526), .B1(n217), .C0(n1513), 
        .C1(n143), .Y(n1188) );
  NAND4X1 U1120 ( .A(n581), .B(n163), .C(n582), .D(n583), .Y(n571) );
  OA21XL U1121 ( .A0(n220), .A1(n587), .B0(n588), .Y(n582) );
  AOI221XL U1122 ( .A0(n76), .A1(n584), .B0(n1664), .B1(n585), .C0(n586), .Y(
        n583) );
  NAND4X1 U1123 ( .A(n932), .B(n152), .C(n933), .D(n934), .Y(n922) );
  OA21XL U1124 ( .A0(n211), .A1(n938), .B0(n939), .Y(n933) );
  AOI221XL U1125 ( .A0(n33), .A1(n142), .B0(n1531), .B1(n144), .C0(n937), .Y(
        n934) );
  NAND4X1 U1126 ( .A(n761), .B(n762), .C(n763), .D(n764), .Y(n757) );
  NAND3X1 U1127 ( .A(n116), .B(n667), .C(n1667), .Y(n763) );
  AOI222XL U1128 ( .A0(n1662), .A1(n155), .B0(n1650), .B1(n253), .C0(n1652), 
        .C1(n1637), .Y(n764) );
  NAND4X1 U1129 ( .A(n1080), .B(n1081), .C(n1082), .D(n1083), .Y(n1076) );
  NAND3X1 U1130 ( .A(n108), .B(n146), .C(n1517), .Y(n1082) );
  AOI222XL U1131 ( .A0(n1514), .A1(n936), .B0(n1536), .B1(n214), .C0(n1518), 
        .C1(n1542), .Y(n1083) );
  NAND4X1 U1132 ( .A(n670), .B(n671), .C(n672), .D(n673), .Y(n659) );
  NAND2X1 U1133 ( .A(n1666), .B(n677), .Y(n670) );
  OAI21XL U1134 ( .A0(n1646), .A1(n1641), .B0(n1659), .Y(n672) );
  AOI222XL U1135 ( .A0(n83), .A1(n674), .B0(n121), .B1(n675), .C0(n676), .C1(
        n180), .Y(n673) );
  NAND4X1 U1136 ( .A(n1021), .B(n1022), .C(n1023), .D(n1024), .Y(n1010) );
  OAI21XL U1137 ( .A0(n1524), .A1(n1537), .B0(n1509), .Y(n1023) );
  NAND2X1 U1138 ( .A(n1502), .B(n1028), .Y(n1021) );
  AOI222XL U1139 ( .A0(n1523), .A1(n1025), .B0(n113), .B1(n1026), .C0(n1027), 
        .C1(n1506), .Y(n1024) );
  NAND4X1 U1140 ( .A(n609), .B(n610), .C(n611), .D(n612), .Y(n605) );
  NAND2X1 U1141 ( .A(n1658), .B(n266), .Y(n611) );
  OAI31XL U1142 ( .A0(n615), .A1(n616), .A2(n617), .B0(n180), .Y(n609) );
  OAI31XL U1143 ( .A0(n1646), .A1(n613), .A2(n614), .B0(n1661), .Y(n610) );
  NAND4X1 U1144 ( .A(n960), .B(n961), .C(n962), .D(n963), .Y(n956) );
  NAND2X1 U1145 ( .A(n1508), .B(n216), .Y(n962) );
  OAI31XL U1146 ( .A0(n966), .A1(n967), .A2(n968), .B0(n165), .Y(n960) );
  OAI31XL U1147 ( .A0(n1524), .A1(n964), .A2(n965), .B0(n1505), .Y(n961) );
  NAND4X1 U1148 ( .A(n788), .B(n598), .C(n789), .D(n790), .Y(n775) );
  NAND3X1 U1149 ( .A(n740), .B(n157), .C(sboxw[26]), .Y(n789) );
  AOI222XL U1150 ( .A0(n1652), .A1(n585), .B0(n1648), .B1(n70), .C0(n76), .C1(
        n74), .Y(n790) );
  NAND4X1 U1151 ( .A(n1107), .B(n949), .C(n1108), .D(n1109), .Y(n1094) );
  NAND3X1 U1152 ( .A(n1059), .B(n1018), .C(sboxw[18]), .Y(n1108) );
  AOI222XL U1153 ( .A0(n1518), .A1(n144), .B0(n1510), .B1(n37), .C0(n33), .C1(
        n35), .Y(n1109) );
  OAI211X1 U1154 ( .A0(n578), .A1(n810), .B0(n811), .C0(n812), .Y(n806) );
  OAI21XL U1155 ( .A0(n613), .A1(n1664), .B0(n1675), .Y(n811) );
  OAI21XL U1156 ( .A0(n813), .A1(n814), .B0(n120), .Y(n812) );
  OAI222XL U1157 ( .A0(n70), .A1(n622), .B0(n154), .B1(n159), .C0(n752), .C1(
        n682), .Y(n814) );
  OAI211X1 U1158 ( .A0(n183), .A1(n1159), .B0(n1160), .C0(n1161), .Y(n1155) );
  OAI21XL U1159 ( .A0(n964), .A1(n1531), .B0(n1506), .Y(n1160) );
  OAI21XL U1160 ( .A0(n1162), .A1(n1163), .B0(n112), .Y(n1161) );
  OAI222XL U1161 ( .A0(n37), .A1(n973), .B0(n143), .B1(n148), .C0(n1071), .C1(
        n1033), .Y(n1163) );
  NAND2X1 U1162 ( .A(n223), .B(n221), .Y(n667) );
  NAND2X1 U1163 ( .A(n266), .B(n221), .Y(n585) );
  NAND2X1 U1164 ( .A(n213), .B(n211), .Y(n1018) );
  NAND2X1 U1165 ( .A(n216), .B(n211), .Y(n936) );
  NAND2X1 U1166 ( .A(n218), .B(n266), .Y(n574) );
  NAND2X1 U1167 ( .A(n208), .B(n216), .Y(n925) );
  NAND2X1 U1168 ( .A(n119), .B(n118), .Y(n600) );
  NAND2X1 U1169 ( .A(n111), .B(n110), .Y(n951) );
  NAND2X1 U1170 ( .A(n82), .B(n117), .Y(n594) );
  NAND2X1 U1171 ( .A(n26), .B(n109), .Y(n945) );
  NAND2X1 U1172 ( .A(n117), .B(n1669), .Y(n753) );
  NAND2X1 U1173 ( .A(n109), .B(n1516), .Y(n1072) );
  NAND2X1 U1174 ( .A(n118), .B(n86), .Y(n645) );
  NAND2X1 U1175 ( .A(n116), .B(n1670), .Y(n622) );
  NAND2X1 U1176 ( .A(n108), .B(n1533), .Y(n973) );
  NAND2X1 U1177 ( .A(n110), .B(n27), .Y(n996) );
  NAND2X1 U1178 ( .A(n102), .B(n100), .Y(n1327) );
  NOR2X1 U1179 ( .A(n657), .B(n266), .Y(n616) );
  NOR2X1 U1180 ( .A(n1008), .B(n216), .Y(n967) );
  NAND2X1 U1181 ( .A(n1663), .B(n221), .Y(n772) );
  NAND2X1 U1182 ( .A(n1522), .B(n211), .Y(n1091) );
  INVX1 U1183 ( .A(n206), .Y(n204) );
  AOI21X1 U1184 ( .A0(n874), .A1(n875), .B0(n858), .Y(n873) );
  AOI222XL U1185 ( .A0(n73), .A1(n1669), .B0(n1662), .B1(n222), .C0(n79), .C1(
        n155), .Y(n874) );
  AOI222XL U1186 ( .A0(n76), .A1(n177), .B0(n219), .B1(n876), .C0(n868), .C1(
        n186), .Y(n875) );
  NAND2X1 U1187 ( .A(n160), .B(n649), .Y(n876) );
  AOI21X1 U1188 ( .A0(n1223), .A1(n1224), .B0(n1207), .Y(n1222) );
  AOI222XL U1189 ( .A0(n39), .A1(n1516), .B0(n1514), .B1(n212), .C0(n30), .C1(
        n936), .Y(n1223) );
  AOI222XL U1190 ( .A0(n33), .A1(n166), .B0(n209), .B1(n1225), .C0(n1217), 
        .C1(n182), .Y(n1224) );
  NAND2X1 U1191 ( .A(n149), .B(n1000), .Y(n1225) );
  OAI222XL U1192 ( .A0(n192), .A1(n297), .B0(n106), .B1(n1378), .C0(n1379), 
        .C1(n168), .Y(n1375) );
  OA21XL U1193 ( .A0(n7), .A1(n5), .B0(n1308), .Y(n1378) );
  OAI22XL U1194 ( .A0(n261), .A1(n205), .B0(n189), .B1(n243), .Y(n1380) );
  NAND2X1 U1195 ( .A(n1337), .B(n203), .Y(n310) );
  NOR4BBX1 U1196 ( .AN(n551), .BN(n397), .C(n558), .D(n559), .Y(n533) );
  OAI2BB2XL U1197 ( .B0(n126), .B1(n375), .A0N(n18), .A1N(n560), .Y(n559) );
  OAI221XL U1198 ( .A0(n201), .A1(n552), .B0(n561), .B1(n173), .C0(n478), .Y(
        n558) );
  AOI211X1 U1199 ( .A0(n1604), .A1(n127), .B0(n562), .C0(n563), .Y(n561) );
  NOR2X1 U1200 ( .A(n244), .B(n205), .Y(n307) );
  INVX1 U1201 ( .A(n227), .Y(n1547) );
  NOR4BX1 U1202 ( .AN(n530), .B(n691), .C(n692), .D(n1618), .Y(n690) );
  OAI21XL U1203 ( .A0(n176), .A1(n403), .B0(n445), .Y(n692) );
  OAI221XL U1204 ( .A0(n21), .A1(n349), .B0(sboxw[1]), .B1(n131), .C0(n693), 
        .Y(n691) );
  AOI222XL U1205 ( .A0(n12), .A1(n136), .B0(n1570), .B1(n205), .C0(n1558), 
        .C1(n191), .Y(n1447) );
  OAI221XL U1206 ( .A0(n177), .A1(n629), .B0(n352), .B1(n575), .C0(n743), .Y(
        n742) );
  OAI221XL U1207 ( .A0(n166), .A1(n980), .B0(n216), .B1(n926), .C0(n1062), .Y(
        n1061) );
  OAI211X1 U1208 ( .A0(n352), .A1(n575), .B0(n815), .C0(n671), .Y(n813) );
  OAI21XL U1209 ( .A0(n76), .A1(n1663), .B0(n186), .Y(n815) );
  OAI211X1 U1210 ( .A0(n217), .A1(n926), .B0(n1164), .C0(n1022), .Y(n1162) );
  OAI21XL U1211 ( .A0(n33), .A1(n1522), .B0(n182), .Y(n1164) );
  AOI211X1 U1212 ( .A0(n1660), .A1(n219), .B0(n889), .C0(n890), .Y(n888) );
  OAI31XL U1213 ( .A0(n624), .A1(n87), .A2(n584), .B0(n661), .Y(n890) );
  OAI222XL U1214 ( .A0(sboxw[25]), .A1(n607), .B0(n121), .B1(n891), .C0(n892), 
        .C1(n180), .Y(n889) );
  AOI211X1 U1215 ( .A0(n1669), .A1(n895), .B0(n616), .C0(n604), .Y(n891) );
  AOI211X1 U1216 ( .A0(n1504), .A1(n209), .B0(n1238), .C0(n1239), .Y(n1237) );
  OAI31XL U1217 ( .A0(n975), .A1(n28), .A2(n142), .B0(n1012), .Y(n1239) );
  OAI222XL U1218 ( .A0(sboxw[17]), .A1(n958), .B0(n113), .B1(n1240), .C0(n1241), .C1(n165), .Y(n1238) );
  AOI211X1 U1219 ( .A0(n1516), .A1(n1244), .B0(n967), .C0(n955), .Y(n1240) );
  OAI211X1 U1220 ( .A0(n737), .A1(n602), .B0(n738), .C0(n739), .Y(n726) );
  AOI32X1 U1221 ( .A0(n740), .A1(n584), .A2(n1666), .B0(n1647), .B1(sboxw[24]), 
        .Y(n739) );
  AOI222XL U1222 ( .A0(n1670), .A1(n158), .B0(n1642), .B1(n81), .C0(n1637), 
        .C1(n83), .Y(n737) );
  OAI21XL U1223 ( .A0(n741), .A1(n742), .B0(n121), .Y(n738) );
  OAI211X1 U1224 ( .A0(n1056), .A1(n953), .B0(n1057), .C0(n1058), .Y(n1045) );
  AOI32X1 U1225 ( .A0(n1059), .A1(n142), .A2(n1502), .B0(n1503), .B1(sboxw[16]), .Y(n1058) );
  AOI222XL U1226 ( .A0(n1533), .A1(n147), .B0(n40), .B1(n32), .C0(n1542), .C1(
        n1523), .Y(n1056) );
  OAI21XL U1227 ( .A0(n1060), .A1(n1061), .B0(n113), .Y(n1057) );
  OAI221XL U1228 ( .A0(n331), .A1(n236), .B0(n106), .B1(n332), .C0(n333), .Y(
        n318) );
  AOI221XL U1229 ( .A0(n48), .A1(n1551), .B0(n1552), .B1(n140), .C0(n335), .Y(
        n333) );
  AOI222XL U1230 ( .A0(n56), .A1(n127), .B0(n1616), .B1(n201), .C0(n1604), 
        .C1(n124), .Y(n699) );
  OAI211X1 U1231 ( .A0(n175), .A1(n349), .B0(n474), .C0(n475), .Y(n470) );
  AOI22X1 U1232 ( .A0(n476), .A1(n174), .B0(n94), .B1(n477), .Y(n475) );
  OAI31XL U1233 ( .A0(n1615), .A1(n1607), .A2(n1626), .B0(n1600), .Y(n474) );
  OAI21XL U1234 ( .A0(n193), .A1(n424), .B0(n131), .Y(n477) );
  NAND2X1 U1235 ( .A(n240), .B(n203), .Y(n1299) );
  OAI222XL U1236 ( .A0(n171), .A1(n244), .B0(sboxw[8]), .B1(n251), .C0(n261), 
        .C1(n191), .Y(n14) );
  OAI221XL U1237 ( .A0(n250), .A1(n267), .B0(n252), .B1(n135), .C0(n268), .Y(
        n265) );
  OAI222XL U1238 ( .A0(n203), .A1(n297), .B0(n106), .B1(n298), .C0(n299), .C1(
        n169), .Y(n293) );
  OAI21XL U1239 ( .A0(n1563), .A1(n303), .B0(n304), .Y(n301) );
  OAI32X1 U1240 ( .A0(n646), .A1(n1642), .A2(n85), .B0(n877), .B1(n663), .Y(
        n872) );
  AOI221XL U1241 ( .A0(n79), .A1(n154), .B0(n73), .B1(n1670), .C0(n878), .Y(
        n877) );
  OAI211X1 U1242 ( .A0(n187), .A1(n159), .B0(n743), .C0(n771), .Y(n878) );
  OAI32X1 U1243 ( .A0(n997), .A1(n40), .A2(n25), .B0(n1226), .B1(n1014), .Y(
        n1221) );
  AOI221XL U1244 ( .A0(n30), .A1(n143), .B0(n39), .B1(n1533), .C0(n1227), .Y(
        n1226) );
  OAI211X1 U1245 ( .A0(n1), .A1(n1072), .B0(n1062), .C0(n1090), .Y(n1227) );
  OAI221XL U1246 ( .A0(n1637), .A1(n87), .B0(sboxw[28]), .B1(sboxw[24]), .C0(
        n118), .Y(n720) );
  OAI221XL U1247 ( .A0(n573), .A1(n222), .B0(n158), .B1(n575), .C0(n576), .Y(
        n572) );
  AOI31X1 U1248 ( .A0(n1642), .A1(n117), .A2(n1667), .B0(n577), .Y(n576) );
  OAI31XL U1249 ( .A0(n186), .A1(n579), .A2(n87), .B0(n580), .Y(n577) );
  OAI221XL U1250 ( .A0(n924), .A1(n212), .B0(n147), .B1(n926), .C0(n927), .Y(
        n923) );
  AOI31X1 U1251 ( .A0(n40), .A1(n109), .A2(n1517), .B0(n928), .Y(n927) );
  OAI31XL U1252 ( .A0(n182), .A1(n930), .A2(n28), .B0(n931), .Y(n928) );
  OAI221XL U1253 ( .A0(n1542), .A1(n28), .B0(n111), .B1(sboxw[16]), .C0(n110), 
        .Y(n1039) );
  AO21X1 U1254 ( .A0(n266), .A1(n1662), .B0(n617), .Y(n675) );
  AO21X1 U1255 ( .A0(n216), .A1(n1514), .B0(n968), .Y(n1026) );
  OAI221XL U1256 ( .A0(n98), .A1(n1326), .B0(n1587), .B1(n1327), .C0(n327), 
        .Y(n1325) );
  OAI221XL U1257 ( .A0(sboxw[28]), .A1(n621), .B0(n622), .B1(n601), .C0(n623), 
        .Y(n619) );
  AOI2BB2X1 U1258 ( .B0(n71), .B1(n1661), .A0N(n70), .A1N(n624), .Y(n621) );
  AOI222XL U1259 ( .A0(n106), .A1(n1353), .B0(n1354), .B1(n168), .C0(n6), .C1(
        n1355), .Y(n1352) );
  NAND4X1 U1260 ( .A(n1293), .B(n1282), .C(n1357), .D(n1358), .Y(n1353) );
  AOI221XL U1261 ( .A0(n1657), .A1(n1642), .B0(n1639), .B1(n637), .C0(n638), 
        .Y(n636) );
  OAI22XL U1262 ( .A0(n120), .A1(n639), .B0(n640), .B1(n1675), .Y(n638) );
  AOI211X1 U1263 ( .A0(n83), .A1(n352), .B0(n641), .C0(n616), .Y(n640) );
  AOI211X1 U1264 ( .A0(n1654), .A1(n186), .B0(n642), .C0(n643), .Y(n639) );
  AOI221XL U1265 ( .A0(n1507), .A1(n40), .B0(n37), .B1(n988), .C0(n989), .Y(
        n987) );
  OAI22XL U1266 ( .A0(n112), .A1(n990), .B0(n991), .B1(n1506), .Y(n989) );
  AOI211X1 U1267 ( .A0(n1523), .A1(n217), .B0(n992), .C0(n967), .Y(n991) );
  AOI211X1 U1268 ( .A0(n1526), .A1(n182), .B0(n993), .C0(n994), .Y(n990) );
  OAI31XL U1269 ( .A0(n1294), .A1(n1295), .A2(n1296), .B0(n1544), .Y(n1267) );
  OAI22XL U1270 ( .A0(n1297), .A1(n236), .B0(n203), .B1(n241), .Y(n1296) );
  OAI211X1 U1271 ( .A0(n201), .A1(n349), .B0(n557), .C0(n445), .Y(n555) );
  OAI21XL U1272 ( .A0(n62), .A1(n1613), .B0(n23), .Y(n557) );
  AOI221XL U1273 ( .A0(n1523), .A1(n212), .B0(n1), .B1(n32), .C0(n1063), .Y(
        n1260) );
  AOI221XL U1274 ( .A0(n1590), .A1(n686), .B0(n1591), .B1(n687), .C0(n688), 
        .Y(n685) );
  NAND4X1 U1275 ( .A(n443), .B(n530), .C(n355), .D(n697), .Y(n687) );
  NAND4X1 U1276 ( .A(n426), .B(n443), .C(n698), .D(n699), .Y(n686) );
  OAI22XL U1277 ( .A0(n689), .A1(n437), .B0(n690), .B1(n409), .Y(n688) );
  OAI31XL U1278 ( .A0(n1649), .A1(sboxw[28]), .A2(n158), .B0(n736), .Y(n799)
         );
  OAI31XL U1279 ( .A0(n574), .A1(sboxw[28]), .A2(n117), .B0(n644), .Y(n643) );
  OAI21XL U1280 ( .A0(n1656), .A1(n79), .B0(n221), .Y(n644) );
  OAI31XL U1281 ( .A0(n925), .A1(n111), .A2(n109), .B0(n995), .Y(n994) );
  OAI21XL U1282 ( .A0(n1513), .A1(n30), .B0(n211), .Y(n995) );
  OAI221XL U1283 ( .A0(n352), .A1(n810), .B0(n819), .B1(n180), .C0(n736), .Y(
        n816) );
  AOI211X1 U1284 ( .A0(n1656), .A1(n157), .B0(n820), .C0(n821), .Y(n819) );
  OAI211X1 U1285 ( .A0(n74), .A1(n573), .B0(n822), .C0(n783), .Y(n820) );
  OAI22XL U1286 ( .A0(n185), .A1(n163), .B0(n70), .B1(n629), .Y(n821) );
  OAI221XL U1287 ( .A0(n217), .A1(n1159), .B0(n1168), .B1(n165), .C0(n1055), 
        .Y(n1165) );
  AOI211X1 U1288 ( .A0(n1513), .A1(n146), .B0(n1169), .C0(n1170), .Y(n1168) );
  OAI211X1 U1289 ( .A0(n35), .A1(n924), .B0(n1171), .C0(n1102), .Y(n1169) );
  OAI22XL U1290 ( .A0(n181), .A1(n926), .B0(n37), .B1(n980), .Y(n1170) );
  AOI211X1 U1291 ( .A0(n76), .A1(n352), .B0(n647), .C0(n648), .Y(n634) );
  OAI22XL U1292 ( .A0(n266), .A1(n649), .B0(n177), .B1(n650), .Y(n648) );
  OAI211X1 U1293 ( .A0(sboxw[24]), .A1(n651), .B0(n652), .C0(n653), .Y(n647)
         );
  AOI211X1 U1294 ( .A0(n33), .A1(n217), .B0(n998), .C0(n999), .Y(n985) );
  OAI22XL U1295 ( .A0(n216), .A1(n1000), .B0(n1542), .B1(n1001), .Y(n999) );
  OAI211X1 U1296 ( .A0(sboxw[16]), .A1(n1002), .B0(n1003), .C0(n1004), .Y(n998) );
  OAI222XL U1297 ( .A0(n765), .A1(n180), .B0(n766), .B1(n747), .C0(n120), .C1(
        n767), .Y(n756) );
  AOI2BB1X1 U1298 ( .A0N(n70), .A1N(n721), .B0(n614), .Y(n766) );
  AOI211X1 U1299 ( .A0(n773), .A1(n219), .B0(n774), .C0(n1664), .Y(n765) );
  AOI211X1 U1300 ( .A0(n1652), .A1(n352), .B0(n768), .C0(n769), .Y(n767) );
  OAI222XL U1301 ( .A0(n1084), .A1(n165), .B0(n1085), .B1(n1066), .C0(n112), 
        .C1(n1086), .Y(n1075) );
  AOI2BB1X1 U1302 ( .A0N(n37), .A1N(n1040), .B0(n965), .Y(n1085) );
  AOI211X1 U1303 ( .A0(n1092), .A1(n209), .B0(n1093), .C0(n1531), .Y(n1084) );
  AOI211X1 U1304 ( .A0(n1518), .A1(n217), .B0(n1087), .C0(n1088), .Y(n1086) );
  OAI211X1 U1305 ( .A0(n911), .A1(n602), .B0(n912), .C0(n913), .Y(n902) );
  AOI2BB2X1 U1306 ( .B0(n914), .B1(n1675), .A0N(n158), .A1N(n628), .Y(n913) );
  AOI32X1 U1307 ( .A0(n121), .A1(n915), .A2(n116), .B0(n1658), .B1(n574), .Y(
        n912) );
  AOI221XL U1308 ( .A0(n83), .A1(n222), .B0(n187), .B1(n81), .C0(n744), .Y(
        n911) );
  AOI32X1 U1309 ( .A0(n113), .A1(n1264), .A2(n108), .B0(n1508), .B1(n925), .Y(
        n1261) );
  OAI21XL U1310 ( .A0(n167), .A1(n1517), .B0(n144), .Y(n1264) );
  OAI211X1 U1311 ( .A0(sboxw[28]), .A1(n154), .B0(n645), .C0(n784), .Y(n781)
         );
  OAI211X1 U1312 ( .A0(n111), .A1(n143), .B0(n996), .C0(n1103), .Y(n1100) );
  AOI211X1 U1313 ( .A0(n1547), .A1(n1444), .B0(n1445), .C0(n1446), .Y(n1443)
         );
  AOI21X1 U1314 ( .A0(n1447), .A1(n1448), .B0(n1313), .Y(n1446) );
  OAI22XL U1315 ( .A0(n1450), .A1(n229), .B0(n1451), .B1(n1315), .Y(n1445) );
  OAI211X1 U1316 ( .A0(n879), .A1(n747), .B0(n880), .C0(n881), .Y(n871) );
  AOI221XL U1317 ( .A0(n80), .A1(n222), .B0(n1669), .B1(n667), .C0(n884), .Y(
        n879) );
  OAI31XL U1318 ( .A0(n615), .A1(n1635), .A2(n730), .B0(n121), .Y(n880) );
  OAI31XL U1319 ( .A0(n882), .A1(n681), .A2(n883), .B0(n180), .Y(n881) );
  OAI211X1 U1320 ( .A0(n1228), .A1(n1066), .B0(n1229), .C0(n1230), .Y(n1220)
         );
  AOI221XL U1321 ( .A0(n31), .A1(n212), .B0(n1516), .B1(n146), .C0(n1233), .Y(
        n1228) );
  OAI31XL U1322 ( .A0(n966), .A1(n1528), .A2(n1049), .B0(n113), .Y(n1229) );
  OAI31XL U1323 ( .A0(n1231), .A1(n1032), .A2(n1232), .B0(n165), .Y(n1230) );
  OAI211X1 U1324 ( .A0(n904), .A1(n180), .B0(n905), .C0(n901), .Y(n903) );
  NAND3X1 U1325 ( .A(n1661), .B(n1668), .C(n178), .Y(n905) );
  NOR4X1 U1326 ( .A(n906), .B(n907), .C(n76), .D(n1636), .Y(n904) );
  OAI221XL U1327 ( .A0(n75), .A1(n628), .B0(n221), .B1(n159), .C0(n908), .Y(
        n906) );
  OAI211X1 U1328 ( .A0(n1253), .A1(n165), .B0(n1254), .C0(n1250), .Y(n1252) );
  NAND3X1 U1329 ( .A(n1505), .B(n1534), .C(n167), .Y(n1254) );
  NOR4X1 U1330 ( .A(n1255), .B(n1256), .C(n33), .D(n1530), .Y(n1253) );
  OAI221XL U1331 ( .A0(n36), .A1(n979), .B0(n211), .B1(n148), .C0(n1257), .Y(
        n1255) );
  OAI211X1 U1332 ( .A0(n594), .A1(n584), .B0(n1633), .C0(n759), .Y(n758) );
  INVX1 U1333 ( .A(n641), .Y(n1633) );
  AOI221XL U1334 ( .A0(n1656), .A1(n75), .B0(n1654), .B1(n1637), .C0(n760), 
        .Y(n759) );
  NOR3X1 U1335 ( .A(n740), .B(n117), .C(n185), .Y(n760) );
  OAI211X1 U1336 ( .A0(n945), .A1(n142), .B0(n1515), .C0(n1078), .Y(n1077) );
  INVX1 U1337 ( .A(n992), .Y(n1515) );
  AOI221XL U1338 ( .A0(n1513), .A1(n36), .B0(n1526), .B1(n1542), .C0(n1079), 
        .Y(n1078) );
  NOR3X1 U1339 ( .A(n1059), .B(sboxw[18]), .C(n181), .Y(n1079) );
  OAI211X1 U1340 ( .A0(n49), .A1(n249), .B0(n1462), .C0(n1339), .Y(n1461) );
  INVX1 U1341 ( .A(n220), .Y(n219) );
  INVX1 U1342 ( .A(n210), .Y(n209) );
  INVX1 U1343 ( .A(n112), .Y(n1506) );
  OAI211X1 U1344 ( .A0(n266), .A1(n160), .B0(n595), .C0(n596), .Y(n593) );
  AND2X2 U1345 ( .A(n597), .B(n598), .Y(n596) );
  OAI211X1 U1346 ( .A0(n215), .A1(n945), .B0(n946), .C0(n947), .Y(n944) );
  AND2X2 U1347 ( .A(n948), .B(n949), .Y(n947) );
  INVX1 U1348 ( .A(n120), .Y(n1675) );
  OAI21XL U1349 ( .A0(sboxw[12]), .A1(n134), .B0(sboxw[11]), .Y(n1346) );
  NAND2X1 U1350 ( .A(n117), .B(sboxw[28]), .Y(n668) );
  NAND2X1 U1351 ( .A(n109), .B(n111), .Y(n1019) );
  OAI21XL U1352 ( .A0(sboxw[28]), .A1(n177), .B0(n118), .Y(n677) );
  OAI21XL U1353 ( .A0(n111), .A1(n1542), .B0(n110), .Y(n1028) );
  OAI22XL U1354 ( .A0(n951), .A1(n211), .B0(n37), .B1(n1040), .Y(n1233) );
  NOR3X1 U1355 ( .A(n602), .B(n1667), .C(n266), .Y(n807) );
  NOR3X1 U1356 ( .A(n953), .B(n1517), .C(n216), .Y(n1156) );
  NAND2X1 U1357 ( .A(n120), .B(n84), .Y(n633) );
  NAND2X1 U1358 ( .A(n112), .B(n25), .Y(n984) );
  NAND2X1 U1359 ( .A(n108), .B(n164), .Y(n975) );
  NAND3X1 U1360 ( .A(n119), .B(n115), .C(n72), .Y(n761) );
  NAND3X1 U1361 ( .A(sboxw[20]), .B(n107), .C(n1541), .Y(n1080) );
  OAI31XL U1362 ( .A0(n657), .A1(n120), .A2(n219), .B0(n603), .Y(n861) );
  OAI31XL U1363 ( .A0(n1008), .A1(n112), .A2(n209), .B0(n954), .Y(n1210) );
  NAND3X1 U1364 ( .A(n482), .B(n127), .C(n89), .Y(n531) );
  NOR2X1 U1365 ( .A(n156), .B(n221), .Y(n744) );
  NOR2X1 U1366 ( .A(n145), .B(n211), .Y(n1063) );
  OAI31XL U1367 ( .A0(n624), .A1(n87), .A2(n220), .B0(n809), .Y(n808) );
  OAI31XL U1368 ( .A0(n975), .A1(n28), .A2(n210), .B0(n1158), .Y(n1157) );
  NOR2X1 U1369 ( .A(n668), .B(n221), .Y(n680) );
  NOR2X1 U1370 ( .A(n1019), .B(n211), .Y(n1031) );
  NAND2X1 U1371 ( .A(n116), .B(n118), .Y(n650) );
  NAND2X1 U1372 ( .A(n108), .B(n110), .Y(n1001) );
  NAND2X1 U1373 ( .A(n1666), .B(n118), .Y(n810) );
  NAND2X1 U1374 ( .A(n1502), .B(n110), .Y(n1159) );
  NOR2X1 U1375 ( .A(n115), .B(n119), .Y(n773) );
  NOR2X1 U1376 ( .A(n107), .B(sboxw[20]), .Y(n1092) );
  INVX1 U1377 ( .A(n260), .Y(n253) );
  INVX1 U1378 ( .A(n215), .Y(n214) );
  INVX1 U1379 ( .A(sboxw[14]), .Y(n42) );
  INVX1 U1380 ( .A(sboxw[30]), .Y(n84) );
  INVX1 U1381 ( .A(sboxw[22]), .Y(n25) );
  OAI221XL U1382 ( .A0(n111), .A1(n972), .B0(n973), .B1(n952), .C0(n974), .Y(
        n970) );
  AOI2BB2X1 U1383 ( .B0(n38), .B1(n1505), .A0N(n37), .A1N(n975), .Y(n972) );
  INVX1 U1384 ( .A(n122), .Y(n85) );
  INVX1 U1385 ( .A(n437), .Y(n1592) );
  INVX1 U1386 ( .A(n663), .Y(n1674) );
  INVX1 U1387 ( .A(n1014), .Y(n1501) );
  INVX1 U1388 ( .A(n858), .Y(n1673) );
  INVX1 U1389 ( .A(n1207), .Y(n1500) );
  NAND2X1 U1390 ( .A(sboxw[14]), .B(n104), .Y(n227) );
  INVX1 U1391 ( .A(n96), .Y(n98) );
  BUFX2 U1392 ( .A(n207), .Y(n206) );
  BUFX2 U1393 ( .A(n207), .Y(n205) );
  INVX1 U1394 ( .A(n104), .Y(n105) );
  INVX1 U1395 ( .A(n99), .Y(n101) );
  NAND2X1 U1396 ( .A(sboxw[14]), .B(sboxw[13]), .Y(n229) );
  BUFX2 U1397 ( .A(sboxw[12]), .Y(n103) );
  AOI222XL U1398 ( .A0(n1485), .A1(n54), .B0(n1591), .B1(n1602), .C0(n95), 
        .C1(n1486), .Y(n1468) );
  AOI211X1 U1399 ( .A0(n1595), .A1(n194), .B0(n1472), .C0(n1473), .Y(n1471) );
  OAI222XL U1400 ( .A0(n406), .A1(n407), .B0(n408), .B1(n409), .C0(n410), .C1(
        n54), .Y(n405) );
  AOI221XL U1401 ( .A0(n432), .A1(n1591), .B0(n433), .B1(n54), .C0(n434), .Y(
        n404) );
  AOI211X1 U1402 ( .A0(n62), .A1(n201), .B0(n421), .C0(n422), .Y(n408) );
  AND2X2 U1403 ( .A(sboxw[0]), .B(n202), .Y(n18) );
  NAND2X1 U1404 ( .A(sboxw[15]), .B(n41), .Y(n1350) );
  INVX1 U1405 ( .A(n104), .Y(n106) );
  BUFX2 U1406 ( .A(n202), .Y(n200) );
  NAND2X1 U1407 ( .A(sboxw[15]), .B(sboxw[14]), .Y(n1266) );
  BUFX2 U1408 ( .A(sboxw[4]), .Y(n92) );
  BUFX2 U1409 ( .A(sboxw[3]), .Y(n91) );
  INVX1 U1410 ( .A(sboxw[15]), .Y(n1543) );
  BUFX2 U1411 ( .A(sboxw[5]), .Y(n93) );
  INVX1 U1412 ( .A(n202), .Y(n198) );
  INVX1 U1413 ( .A(sboxw[0]), .Y(n197) );
  NOR4BX1 U1414 ( .AN(n1278), .B(n1375), .C(n1376), .D(n1557), .Y(n1349) );
  AOI22X1 U1415 ( .A0(sboxw[14]), .A1(n1360), .B0(n1361), .B1(n42), .Y(n1351)
         );
  OAI211X1 U1416 ( .A0(n1370), .A1(n236), .B0(n1371), .C0(n1372), .Y(n1360) );
  NAND2X1 U1417 ( .A(n95), .B(n94), .Y(n437) );
  BUFX2 U1418 ( .A(sboxw[5]), .Y(n94) );
  NAND2X1 U1419 ( .A(n95), .B(n174), .Y(n1113) );
  BUFX2 U1420 ( .A(n202), .Y(n201) );
  INVX1 U1421 ( .A(sboxw[7]), .Y(n1588) );
  AOI222XL U1422 ( .A0(n94), .A1(n460), .B0(n461), .B1(n1597), .C0(n1596), 
        .C1(n462), .Y(n459) );
  AOI221XL U1423 ( .A0(n106), .A1(n1463), .B0(n1464), .B1(n168), .C0(n1465), 
        .Y(n1441) );
  AOI221XL U1424 ( .A0(n94), .A1(n708), .B0(n709), .B1(n1597), .C0(n710), .Y(
        n683) );
  AOI221XL U1425 ( .A0(n74), .A1(n637), .B0(n1671), .B1(n775), .C0(n776), .Y(
        n754) );
  AOI222XL U1426 ( .A0(n122), .A1(n756), .B0(n1671), .B1(n757), .C0(n1672), 
        .C1(n758), .Y(n755) );
  INVX1 U1427 ( .A(n635), .Y(n1671) );
  AOI221XL U1428 ( .A0(n1673), .A1(n658), .B0(n659), .B1(n85), .C0(n660), .Y(
        n630) );
  OAI222XL U1429 ( .A0(n632), .A1(n633), .B0(n634), .B1(n635), .C0(n636), .C1(
        n85), .Y(n631) );
  OAI22XL U1430 ( .A0(n85), .A1(n661), .B0(n662), .B1(n663), .Y(n660) );
  OAI22XL U1431 ( .A0(n122), .A1(n887), .B0(n888), .B1(n85), .Y(n886) );
  AOI222XL U1432 ( .A0(n902), .A1(n85), .B0(n1673), .B1(n1640), .C0(n122), 
        .C1(n903), .Y(n885) );
  AOI211X1 U1433 ( .A0(n1660), .A1(n186), .B0(n896), .C0(n897), .Y(n887) );
  OAI222XL U1434 ( .A0(n857), .A1(n858), .B0(n859), .B1(n663), .C0(n122), .C1(
        n860), .Y(n856) );
  AOI211X1 U1435 ( .A0(n871), .A1(n85), .B0(n872), .C0(n873), .Y(n855) );
  NOR4X1 U1436 ( .A(n861), .B(n862), .C(n863), .D(n864), .Y(n860) );
  OAI22XL U1437 ( .A0(sboxw[23]), .A1(n1073), .B0(n1074), .B1(n374), .Y(
        new_sboxw[20]) );
  AOI221XL U1438 ( .A0(n35), .A1(n988), .B0(n929), .B1(n1094), .C0(n1095), .Y(
        n1073) );
  AOI222XL U1439 ( .A0(n114), .A1(n1075), .B0(n929), .B1(n1076), .C0(n1345), 
        .C1(n1077), .Y(n1074) );
  INVX1 U1440 ( .A(n986), .Y(n929) );
  OAI2BB2XL U1441 ( .B0(sboxw[23]), .B1(n981), .A0N(sboxw[23]), .A1N(n982), 
        .Y(new_sboxw[22]) );
  AOI221XL U1442 ( .A0(n1500), .A1(n1009), .B0(n1010), .B1(n1499), .C0(n1011), 
        .Y(n981) );
  OAI222XL U1443 ( .A0(n983), .A1(n984), .B0(n985), .B1(n986), .C0(n987), .C1(
        n1499), .Y(n982) );
  OAI22XL U1444 ( .A0(n1499), .A1(n1012), .B0(n1013), .B1(n1014), .Y(n1011) );
  OAI2BB2XL U1445 ( .B0(n1204), .B1(n374), .A0N(n1205), .A1N(n374), .Y(
        new_sboxw[17]) );
  OAI222XL U1446 ( .A0(n1206), .A1(n1207), .B0(n1208), .B1(n1014), .C0(n114), 
        .C1(n1209), .Y(n1205) );
  AOI211X1 U1447 ( .A0(n1220), .A1(n1499), .B0(n1221), .C0(n1222), .Y(n1204)
         );
  NOR4X1 U1448 ( .A(n1210), .B(n1211), .C(n1212), .D(n1213), .Y(n1209) );
  OAI2BB2XL U1449 ( .B0(n1234), .B1(n374), .A0N(n1235), .A1N(n374), .Y(
        new_sboxw[16]) );
  AOI222XL U1450 ( .A0(n1251), .A1(n1499), .B0(n1500), .B1(n1511), .C0(n114), 
        .C1(n1252), .Y(n1234) );
  OAI22XL U1451 ( .A0(n114), .A1(n1236), .B0(n1237), .B1(n1499), .Y(n1235) );
  OAI211X1 U1452 ( .A0(n1260), .A1(n953), .B0(n1261), .C0(n1262), .Y(n1251) );
  NOR4BX1 U1453 ( .AN(n841), .B(n842), .C(n843), .D(n1647), .Y(n824) );
  AOI221XL U1454 ( .A0(n121), .A1(n848), .B0(n849), .B1(n1675), .C0(n850), .Y(
        n823) );
  AOI221XL U1455 ( .A0(n1672), .A1(n826), .B0(n1673), .B1(n827), .C0(n828), 
        .Y(n825) );
  NOR3X1 U1456 ( .A(n806), .B(n807), .C(n808), .Y(n792) );
  NOR4BBX1 U1457 ( .AN(n809), .BN(n623), .C(n816), .D(n817), .Y(n791) );
  AOI221XL U1458 ( .A0(n1674), .A1(n794), .B0(n1673), .B1(n795), .C0(n796), 
        .Y(n793) );
  AOI222XL U1459 ( .A0(n121), .A1(n718), .B0(n719), .B1(n1675), .C0(n1661), 
        .C1(n720), .Y(n717) );
  NOR4X1 U1460 ( .A(n745), .B(n746), .C(n1655), .D(n589), .Y(n715) );
  AOI2BB2X1 U1461 ( .B0(n122), .B1(n726), .A0N(n122), .A1N(n727), .Y(n716) );
  AOI211X1 U1462 ( .A0(n120), .A1(n618), .B0(n619), .C0(n620), .Y(n565) );
  AOI211X1 U1463 ( .A0(n604), .A1(n1659), .B0(n605), .C0(n606), .Y(n567) );
  AOI222XL U1464 ( .A0(n570), .A1(n85), .B0(n1674), .B1(n571), .C0(n1673), 
        .C1(n572), .Y(n569) );
  NOR3X1 U1465 ( .A(n548), .B(n549), .C(n550), .Y(n534) );
  NOR4BX1 U1466 ( .AN(n246), .B(n247), .C(n248), .D(n1557), .Y(n228) );
  NOR4X1 U1467 ( .A(n231), .B(n232), .C(n233), .D(n234), .Y(n230) );
  OAI222XL U1468 ( .A0(n1140), .A1(n917), .B0(n1141), .B1(n919), .C0(sboxw[23]), .C1(n1142), .Y(new_sboxw[19]) );
  NOR3X1 U1469 ( .A(n1155), .B(n1156), .C(n1157), .Y(n1141) );
  AOI221XL U1470 ( .A0(n1501), .A1(n1143), .B0(n1500), .B1(n1144), .C0(n1145), 
        .Y(n1142) );
  NOR4BBX1 U1471 ( .AN(n1158), .BN(n974), .C(n1165), .D(n1166), .Y(n1140) );
  OAI222XL U1472 ( .A0(n1172), .A1(n917), .B0(n1173), .B1(n919), .C0(sboxw[23]), .C1(n1174), .Y(new_sboxw[18]) );
  NOR4BX1 U1473 ( .AN(n1190), .B(n1191), .C(n1192), .D(n1503), .Y(n1173) );
  AOI221XL U1474 ( .A0(n113), .A1(n1197), .B0(n1198), .B1(n1506), .C0(n1199), 
        .Y(n1172) );
  AOI221XL U1475 ( .A0(n1345), .A1(n1175), .B0(n1500), .B1(n1176), .C0(n1177), 
        .Y(n1174) );
  AOI211X1 U1476 ( .A0(n112), .A1(n969), .B0(n970), .C0(n971), .Y(n916) );
  AOI211X1 U1477 ( .A0(n955), .A1(n1509), .B0(n956), .C0(n957), .Y(n918) );
  AOI222XL U1478 ( .A0(n921), .A1(n1499), .B0(n1501), .B1(n922), .C0(n1500), 
        .C1(n923), .Y(n920) );
  OAI222XL U1479 ( .A0(n1034), .A1(n919), .B0(sboxw[23]), .B1(n1035), .C0(
        n1036), .C1(n917), .Y(new_sboxw[21]) );
  AOI222XL U1480 ( .A0(n113), .A1(n1037), .B0(n1038), .B1(n1506), .C0(n1505), 
        .C1(n1039), .Y(n1036) );
  NOR4X1 U1481 ( .A(n1064), .B(n1065), .C(n1512), .D(n940), .Y(n1034) );
  AOI2BB2X1 U1482 ( .B0(n114), .B1(n1045), .A0N(n114), .A1N(n1046), .Y(n1035)
         );
  AOI222XL U1483 ( .A0(n95), .A1(n498), .B0(n1589), .B1(n499), .C0(n1590), 
        .C1(n500), .Y(n497) );
  AOI222XL U1484 ( .A0(sboxw[14]), .A1(n1383), .B0(n1546), .B1(n1384), .C0(
        n1545), .C1(n1385), .Y(n1382) );
  AOI221XL U1485 ( .A0(n1547), .A1(n1330), .B0(n1331), .B1(n42), .C0(n1332), 
        .Y(n1310) );
  AOI222XL U1486 ( .A0(n318), .A1(n42), .B0(n1547), .B1(n1556), .C0(sboxw[14]), 
        .C1(n319), .Y(n289) );
  OAI22XL U1487 ( .A0(sboxw[14]), .A1(n291), .B0(n292), .B1(n42), .Y(n290) );
  AOI211X1 U1488 ( .A0(n1550), .A1(sboxw[8]), .B0(n293), .C0(n294), .Y(n292)
         );
  AOI211X1 U1489 ( .A0(n1550), .A1(n50), .B0(n308), .C0(n309), .Y(n291) );
  OAI31XL U1490 ( .A0(n295), .A1(n45), .A2(n4), .B0(n296), .Y(n294) );
  BUFX2 U1491 ( .A(n222), .Y(n220) );
  BUFX2 U1492 ( .A(n352), .Y(n260) );
  BUFX2 U1493 ( .A(n212), .Y(n210) );
  BUFX2 U1494 ( .A(n217), .Y(n215) );
  BUFX2 U1495 ( .A(n222), .Y(n221) );
  BUFX2 U1496 ( .A(n212), .Y(n211) );
  BUFX2 U1497 ( .A(n352), .Y(n266) );
  BUFX2 U1498 ( .A(n217), .Y(n216) );
  BUFX2 U1499 ( .A(sboxw[19]), .Y(n110) );
  BUFX2 U1500 ( .A(sboxw[27]), .Y(n118) );
  AOI2BB2X1 U1501 ( .B0(n95), .B1(n468), .A0N(n95), .A1N(n469), .Y(n458) );
  NOR4X1 U1502 ( .A(n470), .B(n471), .C(n472), .D(n1611), .Y(n469) );
  BUFX2 U1503 ( .A(sboxw[21]), .Y(n112) );
  BUFX2 U1504 ( .A(sboxw[29]), .Y(n120) );
  BUFX2 U1505 ( .A(sboxw[28]), .Y(n119) );
  BUFX2 U1506 ( .A(sboxw[20]), .Y(n111) );
  OAI222XL U1507 ( .A0(n1112), .A1(n1113), .B0(n1114), .B1(n437), .C0(n95), 
        .C1(n1115), .Y(n1111) );
  NOR4X1 U1508 ( .A(n1124), .B(n1125), .C(n391), .D(n1611), .Y(n1112) );
  NOR4X1 U1509 ( .A(n1116), .B(n1117), .C(n1118), .D(n1119), .Y(n1115) );
  NOR4BX1 U1510 ( .AN(n514), .B(n1121), .C(n1122), .D(n1603), .Y(n1114) );
  AOI211X1 U1511 ( .A0(n1629), .A1(n59), .B0(n493), .C0(n1612), .Y(n492) );
  OAI22XL U1512 ( .A0(n202), .A1(n126), .B0(n1629), .B1(n131), .Y(n493) );
  INVX1 U1513 ( .A(n485), .Y(n1612) );
  NAND2X1 U1514 ( .A(n122), .B(n121), .Y(n663) );
  NAND2X1 U1515 ( .A(n114), .B(n113), .Y(n1014) );
  NAND2X1 U1516 ( .A(n122), .B(n179), .Y(n858) );
  NAND2X1 U1517 ( .A(n114), .B(n164), .Y(n1207) );
  INVX1 U1518 ( .A(n114), .Y(n1499) );
  BUFX2 U1519 ( .A(sboxw[21]), .Y(n113) );
  BUFX2 U1520 ( .A(sboxw[29]), .Y(n121) );
  NAND2X1 U1521 ( .A(n95), .B(sboxw[7]), .Y(n340) );
  NAND2X1 U1522 ( .A(sboxw[7]), .B(n53), .Y(n342) );
  NAND2X1 U1523 ( .A(sboxw[31]), .B(n84), .Y(n568) );
  NAND2X1 U1524 ( .A(sboxw[23]), .B(n25), .Y(n919) );
  NAND2X1 U1525 ( .A(n122), .B(sboxw[31]), .Y(n566) );
  NAND2X1 U1526 ( .A(n114), .B(sboxw[23]), .Y(n917) );
  INVX1 U1527 ( .A(sboxw[31]), .Y(n1631) );
  INVX1 U1528 ( .A(sboxw[23]), .Y(n374) );
  INVX1 U1529 ( .A(sboxw[13]), .Y(n104) );
  BUFX2 U1530 ( .A(sboxw[6]), .Y(n95) );
  INVX1 U1531 ( .A(sboxw[24]), .Y(n222) );
  INVX1 U1532 ( .A(sboxw[25]), .Y(n352) );
  INVX1 U1533 ( .A(sboxw[16]), .Y(n212) );
  INVX1 U1534 ( .A(sboxw[17]), .Y(n217) );
  BUFX2 U1535 ( .A(sboxw[30]), .Y(n122) );
  BUFX2 U1536 ( .A(sboxw[22]), .Y(n114) );
  OAI211X1 U1537 ( .A0(n1265), .A1(n1266), .B0(n1267), .C0(n1268), .Y(
        new_sboxw[15]) );
  OAI222XL U1538 ( .A0(n683), .A1(n340), .B0(n684), .B1(n342), .C0(sboxw[7]), 
        .C1(n685), .Y(new_sboxw[2]) );
  OAI222XL U1539 ( .A0(n533), .A1(n340), .B0(n534), .B1(n342), .C0(sboxw[7]), 
        .C1(n535), .Y(new_sboxw[3]) );
  OAI222XL U1540 ( .A0(n457), .A1(n342), .B0(sboxw[7]), .B1(n458), .C0(n459), 
        .C1(n340), .Y(new_sboxw[5]) );
  OAI222XL U1541 ( .A0(n1349), .A1(n1350), .B0(sboxw[15]), .B1(n1351), .C0(
        n1352), .C1(n1266), .Y(new_sboxw[13]) );
  OAI222XL U1542 ( .A0(n1441), .A1(n1266), .B0(n1442), .B1(n1350), .C0(
        sboxw[15]), .C1(n1443), .Y(new_sboxw[10]) );
  OAI222XL U1543 ( .A0(n339), .A1(n340), .B0(n341), .B1(n342), .C0(sboxw[7]), 
        .C1(n343), .Y(new_sboxw[7]) );
  OAI2BB2XL U1544 ( .B0(n289), .B1(n1543), .A0N(n290), .A1N(n1543), .Y(
        new_sboxw[8]) );
  OAI22XL U1545 ( .A0(sboxw[7]), .A1(n496), .B0(n497), .B1(n1588), .Y(
        new_sboxw[4]) );
  OAI2BB2XL U1546 ( .B0(n1110), .B1(n1588), .A0N(n1111), .A1N(n1588), .Y(
        new_sboxw[1]) );
  OAI2BB2XL U1547 ( .B0(sboxw[15]), .B1(n1310), .A0N(sboxw[15]), .A1N(n1311), 
        .Y(new_sboxw[14]) );
  OAI22XL U1548 ( .A0(n1381), .A1(sboxw[15]), .B0(n1382), .B1(n1543), .Y(
        new_sboxw[12]) );
  OAI2BB2XL U1549 ( .B0(n224), .B1(n1543), .A0N(n225), .A1N(n1543), .Y(
        new_sboxw[9]) );
  OAI2BB1X1 U1550 ( .A0N(n1327), .A1N(n287), .B0(n191), .Y(n1406) );
  AOI221XL U1551 ( .A0(n44), .A1(n51), .B0(n46), .B1(n141), .C0(n338), .Y(n331) );
  AOI222XL U1552 ( .A0(n170), .A1(n44), .B0(n172), .B1(n1359), .C0(n190), .C1(
        n1558), .Y(n1358) );
  AOI221XL U1553 ( .A0(n13), .A1(n1562), .B0(n44), .B1(n192), .C0(n1402), .Y(
        n1401) );
  NAND3XL U1554 ( .A(n44), .B(n191), .C(n1553), .Y(n1278) );
  NAND4BX1 U1555 ( .AN(n454), .B(n503), .C(n17), .D(n545), .Y(n537) );
  NAND4X1 U1556 ( .A(n513), .B(n371), .C(n514), .D(n504), .Y(n510) );
  AOI21XL U1557 ( .A0(n125), .A1(n56), .B0(n388), .Y(n508) );
  AOI211XL U1558 ( .A0(n1334), .A1(n45), .B0(n1335), .C0(n328), .Y(n1333) );
  NAND2X1 U1559 ( .A(n1579), .B(n52), .Y(n1282) );
  OAI2BB2XL U1560 ( .B0(n203), .B1(n281), .A0N(n134), .A1N(n1581), .Y(n280) );
  AOI222XL U1561 ( .A0(n48), .A1(n1574), .B0(n1554), .B1(n1586), .C0(n1564), 
        .C1(n5), .Y(n1410) );
  INVX1 U1562 ( .A(n1281), .Y(n1559) );
  OAI211XL U1563 ( .A0(n50), .A1(n288), .B0(n1356), .C0(n1281), .Y(n1354) );
  NAND2XL U1564 ( .A(n288), .B(n281), .Y(n1467) );
  NOR2XL U1565 ( .A(n281), .B(n96), .Y(n1347) );
  NAND3X1 U1566 ( .A(n1596), .B(n1623), .C(n176), .Y(n1488) );
  OAI2BB2XL U1567 ( .B0(n22), .B1(n19), .A0N(n1623), .A1N(n128), .Y(n450) );
  NAND3X1 U1568 ( .A(n20), .B(n1623), .C(n1593), .Y(n364) );
  OAI21XL U1569 ( .A0(n65), .A1(n1623), .B0(n123), .Y(n473) );
  NAND2X1 U1570 ( .A(n63), .B(n1623), .Y(n361) );
  NAND3XL U1571 ( .A(n100), .B(n135), .C(n1563), .Y(n1390) );
  AOI211XL U1572 ( .A0(n49), .A1(n100), .B0(n1418), .C0(n1419), .Y(n1417) );
  NAND3XL U1573 ( .A(n337), .B(n135), .C(n100), .Y(n1409) );
  OAI21XL U1574 ( .A0(n97), .A1(n1327), .B0(n133), .Y(n1365) );
  OAI221XL U1575 ( .A0(n172), .A1(n139), .B0(n204), .B1(n133), .C0(n1454), .Y(
        n1452) );
  OAI222XL U1576 ( .A0(n171), .A1(n139), .B0(n50), .B1(n316), .C0(n136), .C1(
        n133), .Y(n1440) );
  AOI211XL U1577 ( .A0(n1555), .A1(n98), .B0(n1397), .C0(n1579), .Y(n1392) );
  NOR2XL U1578 ( .A(n330), .B(n1579), .Y(n1431) );
  AOI221XL U1579 ( .A0(n98), .A1(n1566), .B0(n1579), .B1(n171), .C0(n1426), 
        .Y(n1421) );
  AOI21X1 U1580 ( .A0(n1129), .A1(n1130), .B0(n1113), .Y(n1128) );
  OAI32X1 U1581 ( .A0(n420), .A1(n1629), .A2(n54), .B0(n1132), .B1(n437), .Y(
        n1127) );
  OAI222XL U1582 ( .A0(n98), .A1(n252), .B0(n283), .B1(n96), .C0(n50), .C1(
        n244), .Y(n1418) );
  OAI21XL U1583 ( .A0(n283), .A1(n4), .B0(n317), .Y(n1424) );
  NOR3X1 U1584 ( .A(n337), .B(n101), .C(n13), .Y(n1387) );
  OAI22XL U1585 ( .A0(n1416), .A1(n227), .B0(n1417), .B1(n229), .Y(n1415) );
  OAI222XL U1586 ( .A0(n226), .A1(n227), .B0(n228), .B1(n229), .C0(sboxw[14]), 
        .C1(n230), .Y(n225) );
  AND2X2 U1587 ( .A(n358), .B(n125), .Y(n15) );
  NAND4X1 U1588 ( .A(n327), .B(n281), .C(n1406), .D(n1407), .Y(n1403) );
  OAI22XL U1589 ( .A0(n139), .A1(n141), .B0(n96), .B1(n316), .Y(n1425) );
  OAI22XL U1590 ( .A0(n334), .A1(n316), .B0(n1289), .B1(n52), .Y(n1284) );
  OAI221XL U1591 ( .A0(n206), .A1(n316), .B0(n172), .B1(n139), .C0(n272), .Y(
        n1374) );
  NAND2X1 U1592 ( .A(n1337), .B(n135), .Y(n296) );
  OAI211X1 U1593 ( .A0(n1134), .A1(n489), .B0(n1135), .C0(n1136), .Y(n1126) );
  BUFX2 U1594 ( .A(n267), .Y(n141) );
  AOI211X1 U1595 ( .A0(n278), .A1(n101), .B0(n279), .C0(n280), .Y(n277) );
  NAND2X1 U1596 ( .A(n560), .B(n127), .Y(n435) );
  AOI211XL U1597 ( .A0(n190), .A1(n1573), .B0(n1380), .C0(n1565), .Y(n1379) );
  NAND2X1 U1598 ( .A(n13), .B(n1573), .Y(n1368) );
  AOI2BB2X1 U1599 ( .B0(n1573), .B1(sboxw[8]), .A0N(n243), .A1N(n190), .Y(n242) );
  AOI221XL U1600 ( .A0(n134), .A1(n1580), .B0(n1562), .B1(n192), .C0(n1571), 
        .Y(n1300) );
  AOI211XL U1601 ( .A0(n1580), .A1(n1321), .B0(n1322), .C0(n1323), .Y(n1318)
         );
  NOR4BXL U1602 ( .AN(n1388), .B(n1420), .C(n1347), .D(n1580), .Y(n1416) );
  NAND4BXL U1603 ( .AN(n1292), .B(n1336), .C(n1408), .D(n1457), .Y(n1444) );
  OAI211XL U1604 ( .A0(sboxw[9]), .A1(n244), .B0(n1336), .C0(n1454), .Y(n1463)
         );
  INVX1 U1605 ( .A(n1336), .Y(n1578) );
  NAND2X1 U1606 ( .A(n1579), .B(sboxw[8]), .Y(n1336) );
  NOR2X1 U1607 ( .A(n63), .B(n92), .Y(n515) );
  NAND3XL U1608 ( .A(n92), .B(n63), .C(n68), .Y(n503) );
  NAND2X1 U1609 ( .A(n1593), .B(n451), .Y(n444) );
  NAND2X1 U1610 ( .A(sboxw[3]), .B(n63), .Y(n512) );
  BUFX2 U1611 ( .A(n17), .Y(n19) );
  NOR4XL U1612 ( .A(n300), .B(n301), .C(n43), .D(n1575), .Y(n299) );
  AOI221XL U1613 ( .A0(n1586), .A1(n12), .B0(n1562), .B1(n306), .C0(n307), .Y(
        n298) );
  AOI222XL U1614 ( .A0(n1580), .A1(n334), .B0(n190), .B1(n46), .C0(n172), .C1(
        n44), .Y(n1370) );
  AOI211X1 U1615 ( .A0(n12), .A1(n206), .B0(n1320), .C0(n307), .Y(n1319) );
  INVXL U1616 ( .A(n1320), .Y(n1561) );
  OAI211X1 U1617 ( .A0(n284), .A1(n192), .B0(n1561), .C0(n1386), .Y(n1385) );
  AOI221XL U1618 ( .A0(n48), .A1(n1558), .B0(n1587), .B1(n1570), .C0(n1387), 
        .Y(n1386) );
  NAND4BX1 U1619 ( .AN(n378), .B(n372), .C(n362), .D(n465), .Y(n460) );
  INVX1 U1620 ( .A(n362), .Y(n1617) );
  OAI211X1 U1621 ( .A0(n201), .A1(n424), .B0(n362), .C0(n495), .Y(n521) );
  INVX1 U1622 ( .A(n15), .Y(n20) );
  OAI31XL U1623 ( .A0(n275), .A1(sboxw[11]), .A2(n5), .B0(n1299), .Y(n1295) );
  AOI211X1 U1624 ( .A0(n1609), .A1(n201), .B0(n510), .C0(n511), .Y(n509) );
  OAI32X1 U1625 ( .A0(n269), .A1(n190), .A2(n42), .B0(n270), .B1(n229), .Y(
        n263) );
  OAI211X1 U1626 ( .A0(n1494), .A1(n376), .B0(n1495), .C0(n1496), .Y(n1485) );
  NOR4X1 U1627 ( .A(n1489), .B(n1490), .C(n62), .D(n11), .Y(n1487) );
  OAI31XL U1628 ( .A0(n398), .A1(n58), .A2(n123), .B0(n435), .Y(n1473) );
  NAND4X1 U1629 ( .A(n1408), .B(n1282), .C(n1409), .D(n1410), .Y(n1398) );
  NOR3XL U1630 ( .A(n1568), .B(n50), .C(n1288), .Y(n1285) );
  AOI2BB2XL U1631 ( .B0(n1497), .B1(n174), .A0N(n348), .A1N(n402), .Y(n1496)
         );
  AOI32XL U1632 ( .A0(n94), .A1(n1498), .A2(n90), .B0(n1599), .B1(n128), .Y(
        n1495) );
  AOI211XL U1633 ( .A0(n22), .A1(n61), .B0(n542), .C0(n543), .Y(n539) );
  AOI32XL U1634 ( .A0(n7), .A1(n47), .A2(n172), .B0(n323), .B1(n49), .Y(n1457)
         );
  AO22X1 U1635 ( .A0(n101), .A1(n278), .B0(n267), .B1(n323), .Y(n1449) );
  AOI211XL U1636 ( .A0(n323), .A1(n1586), .B0(n324), .C0(n325), .Y(n320) );
  NOR2X1 U1637 ( .A(n126), .B(n198), .Y(n388) );
  AOI211X1 U1638 ( .A0(n93), .A1(n392), .B0(n393), .C0(n394), .Y(n339) );
  NOR3X1 U1639 ( .A(n376), .B(n60), .C(n176), .Y(n703) );
  NOR3X1 U1640 ( .A(n376), .B(n1608), .C(n200), .Y(n549) );
  OAI211X1 U1641 ( .A0(n479), .A1(n376), .B0(n480), .C0(n481), .Y(n468) );
  OAI21XL U1642 ( .A0(n58), .A1(n376), .B0(n377), .Y(n373) );
  NAND2XL U1643 ( .A(n560), .B(n198), .Y(n701) );
  NOR2XL U1644 ( .A(n376), .B(n494), .Y(n560) );
  AOI221XL U1645 ( .A0(n59), .A1(n124), .B0(n69), .B1(n8), .C0(n1133), .Y(
        n1132) );
  OAI31XL U1646 ( .A0(n1137), .A1(n455), .A2(n1138), .B0(n173), .Y(n1136) );
  OAI2BB1X1 U1647 ( .A0N(n58), .A1N(n127), .B0(n91), .Y(n451) );
  NAND3X1 U1648 ( .A(n1583), .B(n191), .C(n103), .Y(n1462) );
  NOR4BXL U1649 ( .AN(n1476), .B(n1477), .C(n1613), .D(n472), .Y(n1475) );
  OAI21XL U1650 ( .A0(n1604), .A1(n59), .B0(n195), .Y(n418) );
  NOR2X1 U1651 ( .A(n442), .B(n195), .Y(n454) );
  NOR2X1 U1652 ( .A(n126), .B(n195), .Y(n486) );
  AOI22XL U1653 ( .A0(n24), .A1(n529), .B0(n1626), .B1(n90), .Y(n698) );
  NAND2X1 U1654 ( .A(n529), .B(n193), .Y(n696) );
  INVXL U1655 ( .A(n415), .Y(n1606) );
  AOI211XL U1656 ( .A0(n56), .A1(n201), .B0(n415), .C0(n390), .Y(n414) );
  AOI221XL U1657 ( .A0(n56), .A1(n196), .B0(n15), .B1(n61), .C0(n486), .Y(
        n1494) );
  AOI221XL U1658 ( .A0(n1573), .A1(n48), .B0(n306), .B1(n1562), .C0(n330), .Y(
        n329) );
  OAI211X1 U1659 ( .A0(n206), .A1(n1327), .B0(n1293), .C0(n138), .Y(n1402) );
  AOI221XL U1660 ( .A0(n43), .A1(n135), .B0(n1560), .B1(n10), .C0(n1576), .Y(
        n332) );
  OAI2BB1X1 U1661 ( .A0N(n10), .A1N(n326), .B0(n327), .Y(n325) );
  AOI211X1 U1662 ( .A0(n336), .A1(n10), .B0(n99), .C0(n168), .Y(n335) );
  AOI211X1 U1663 ( .A0(n42), .A1(n262), .B0(n264), .C0(n263), .Y(n224) );
  OAI2BB2XL U1664 ( .B0(n261), .B1(n1276), .A0N(n1585), .A1N(n1337), .Y(n1437)
         );
  OAI21XL U1665 ( .A0(n48), .A1(n261), .B0(n1368), .Y(n1364) );
  AOI32XL U1666 ( .A0(n337), .A1(n192), .A2(n1549), .B0(n1548), .B1(sboxw[8]), 
        .Y(n1372) );
  OAI211XL U1667 ( .A0(sboxw[12]), .A1(n192), .B0(n261), .C0(n235), .Y(n1404)
         );
  OAI222XL U1668 ( .A0(n5), .A1(n133), .B0(sboxw[8]), .B1(n251), .C0(n7), .C1(
        n1342), .Y(n1423) );
  OAI222XL U1669 ( .A0(n171), .A1(n133), .B0(n251), .B1(n192), .C0(n7), .C1(
        n1321), .Y(n1433) );
  OAI221XL U1670 ( .A0(sboxw[12]), .A1(n1305), .B0(n133), .B1(n1276), .C0(
        n1306), .Y(n1303) );
  OAI31XL U1671 ( .A0(n1583), .A1(sboxw[12]), .A2(n334), .B0(n1368), .Y(n1426)
         );
  OAI31XL U1672 ( .A0(n1583), .A1(sboxw[12]), .A2(n1586), .B0(n1408), .Y(n1419) );
  OAI221XL U1673 ( .A0(n1587), .A1(n45), .B0(n98), .B1(sboxw[12]), .C0(
        sboxw[11]), .Y(n1355) );
  AOI211X1 U1674 ( .A0(n1564), .A1(n206), .B0(n1395), .C0(n1396), .Y(n1394) );
  OAI222XL U1675 ( .A0(n1312), .A1(n1313), .B0(n1314), .B1(n1315), .C0(n1316), 
        .C1(n42), .Y(n1311) );
  AOI32XL U1676 ( .A0(n494), .A1(n64), .A2(n1630), .B0(n529), .B1(n18), .Y(
        n697) );
  OA21XL U1677 ( .A0(n494), .A1(n359), .B0(n400), .Y(n491) );
  NAND4X1 U1678 ( .A(n503), .B(n504), .C(n505), .D(n506), .Y(n499) );
  OAI221XL U1679 ( .A0(n92), .A1(n395), .B0(n131), .B1(n375), .C0(n397), .Y(
        n393) );
  OAI221XL U1680 ( .A0(n1630), .A1(n58), .B0(sboxw[4]), .B1(sboxw[0]), .C0(n91), .Y(n462) );
  OAI31XL U1681 ( .A0(n1624), .A1(sboxw[4]), .A2(n348), .B0(n478), .Y(n541) );
  OAI32XL U1682 ( .A0(n196), .A1(sboxw[4]), .A2(n90), .B0(n69), .B1(n512), .Y(
        n1125) );
  OAI31XL U1683 ( .A0(n128), .A1(sboxw[4]), .A2(sboxw[2]), .B0(n418), .Y(n417)
         );
  OAI211X1 U1684 ( .A0(sboxw[4]), .A1(n124), .B0(n126), .C0(n526), .Y(n523) );
  OAI222XL U1685 ( .A0(n1300), .A1(n169), .B0(sboxw[13]), .B1(n1301), .C0(n141), .C1(n297), .Y(n1294) );
  OAI31XL U1686 ( .A0(n295), .A1(sboxw[11]), .A2(n141), .B0(n1278), .Y(n1274)
         );
  OAI22XL U1687 ( .A0(n95), .A1(n1470), .B0(n1471), .B1(n54), .Y(n1469) );
  NAND2X1 U1688 ( .A(n198), .B(n411), .Y(n386) );
  OAI211XL U1689 ( .A0(sboxw[1]), .A1(n431), .B0(n443), .C0(n693), .Y(n708) );
  OAI211X1 U1690 ( .A0(n67), .A1(n431), .B0(n514), .C0(n525), .Y(n524) );
  AOI2BB2X1 U1691 ( .B0(n91), .B1(n199), .A0N(n199), .A1N(n494), .Y(n526) );
  OAI211X1 U1692 ( .A0(n20), .A1(n463), .B0(n464), .C0(n371), .Y(n461) );
  OAI221XL U1693 ( .A0(n175), .A1(n403), .B0(n201), .B1(n349), .C0(n485), .Y(
        n484) );
  OAI211X1 U1694 ( .A0(n15), .A1(n495), .B0(n485), .C0(n513), .Y(n1133) );
  AOI222XL U1695 ( .A0(n8), .A1(n348), .B0(n1629), .B1(n61), .C0(n1630), .C1(
        n56), .Y(n479) );
  AOI222XL U1696 ( .A0(n68), .A1(n1620), .B0(n175), .B1(n515), .C0(n194), .C1(
        n56), .Y(n1476) );
  AOI221XL U1697 ( .A0(n60), .A1(n196), .B0(n1607), .B1(n441), .C0(n1139), .Y(
        n1134) );
  AOI222XL U1698 ( .A0(n1586), .A1(n46), .B0(n323), .B1(n134), .C0(n98), .C1(
        n1558), .Y(n1407) );
  OAI211X1 U1699 ( .A0(n1627), .A1(n126), .B0(n1622), .C0(n452), .Y(n432) );
  OAI222XL U1700 ( .A0(n126), .A1(n16), .B0(n130), .B1(n123), .C0(n1627), .C1(
        n19), .Y(n416) );
  INVX1 U1701 ( .A(n456), .Y(n1627) );
  AOI2BB2X1 U1702 ( .B0(n1609), .B1(n193), .A0N(n123), .A1N(n402), .Y(n544) );
  XOR2X1 U1703 ( .A(n64), .B(n193), .Y(n1493) );
  OAI222XL U1704 ( .A0(n258), .A1(n140), .B0(n98), .B1(n305), .C0(n288), .C1(
        n1342), .Y(n1420) );
  NAND4BX1 U1705 ( .AN(n315), .B(n1282), .C(n284), .D(n1466), .Y(n1464) );
  OAI21XL U1706 ( .A0(n170), .A1(n284), .B0(n1282), .Y(n1307) );
  AOI2BB2X1 U1707 ( .B0(n43), .B1(n204), .A0N(n172), .A1N(n138), .Y(n1454) );
endmodule


module aes_core ( clk, reset_n, encdec, init, next, ready, key, keylen, block, 
        result, result_valid );
  input [255:0] key;
  input [127:0] block;
  output [127:0] result;
  input clk, reset_n, encdec, init, next, keylen;
  output ready, result_valid;
  wire   enc_next, enc_ready, dec_next, dec_ready, key_ready, n4, n5, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n1, n2, n3, n6,
         n7, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83;
  wire   [3:0] enc_round_nr;
  wire   [127:0] round_key;
  wire   [31:0] enc_sboxw;
  wire   [31:0] new_sboxw;
  wire   [127:0] enc_new_block;
  wire   [3:0] dec_round_nr;
  wire   [127:0] dec_new_block;
  wire   [3:0] muxed_round_nr;
  wire   [31:0] keymem_sboxw;
  wire   [31:0] muxed_sboxw;
  wire   [1:0] aes_core_ctrl_reg;

  aes_encipher_block enc_block ( .clk(clk), .reset_n(n80), .next(enc_next), 
        .keylen(keylen), .round(enc_round_nr), .round_key(round_key), .sboxw(
        enc_sboxw), .new_sboxw({new_sboxw[31:16], n3, n38, n26, n40, n1, n28, 
        n42, n32, n30, new_sboxw[6], n24, n34, n22, n7, n36, new_sboxw[0]}), 
        .block(block), .new_block(enc_new_block), .ready(enc_ready) );
  aes_decipher_block dec_block ( .clk(clk), .reset_n(n80), .next(dec_next), 
        .keylen(keylen), .round(dec_round_nr), .round_key(round_key), .block(
        block), .new_block(dec_new_block), .ready(dec_ready) );
  aes_key_mem keymem ( .clk(clk), .reset_n(n80), .key(key), .keylen(keylen), 
        .init(init), .round(muxed_round_nr), .round_key(round_key), .ready(
        key_ready), .sboxw(keymem_sboxw), .new_sboxw(new_sboxw) );
  aes_sbox sbox_inst ( .sboxw(muxed_sboxw), .new_sboxw(new_sboxw) );
  DFFRX1 result_valid_reg_reg ( .D(n17), .CK(clk), .RN(n80), .Q(result_valid)
         );
  DFFSX1 ready_reg_reg ( .D(n18), .CK(clk), .SN(n80), .Q(ready) );
  DFFRX1 \aes_core_ctrl_reg_reg[1]  ( .D(n19), .CK(clk), .RN(n80), .Q(
        aes_core_ctrl_reg[1]), .QN(n4) );
  DFFRX1 \aes_core_ctrl_reg_reg[0]  ( .D(n20), .CK(clk), .RN(n80), .Q(
        aes_core_ctrl_reg[0]), .QN(n5) );
  BUFX2 U3 ( .A(reset_n), .Y(n80) );
  AO22X1 U4 ( .A0(keymem_sboxw[11]), .A1(n44), .B0(enc_sboxw[11]), .B1(n47), 
        .Y(muxed_sboxw[11]) );
  AO22X1 U5 ( .A0(keymem_sboxw[12]), .A1(n44), .B0(enc_sboxw[12]), .B1(n47), 
        .Y(muxed_sboxw[12]) );
  AO22X1 U6 ( .A0(keymem_sboxw[8]), .A1(n43), .B0(n48), .B1(enc_sboxw[8]), .Y(
        muxed_sboxw[8]) );
  AO22X1 U7 ( .A0(keymem_sboxw[9]), .A1(n43), .B0(n48), .B1(enc_sboxw[9]), .Y(
        muxed_sboxw[9]) );
  INVX1 U8 ( .A(n33), .Y(n34) );
  INVX1 U9 ( .A(n39), .Y(n40) );
  INVX1 U10 ( .A(n2), .Y(n3) );
  INVX1 U11 ( .A(n6), .Y(n7) );
  INVX1 U12 ( .A(n31), .Y(n32) );
  INVX1 U13 ( .A(n27), .Y(n28) );
  INVX1 U14 ( .A(n23), .Y(n24) );
  INVX1 U15 ( .A(n35), .Y(n36) );
  INVX1 U16 ( .A(n41), .Y(n42) );
  INVX1 U17 ( .A(n25), .Y(n26) );
  INVX1 U18 ( .A(n21), .Y(n22) );
  BUFX2 U19 ( .A(new_sboxw[11]), .Y(n1) );
  INVX1 U20 ( .A(n37), .Y(n38) );
  INVX1 U21 ( .A(n29), .Y(n30) );
  AO22X1 U22 ( .A0(keymem_sboxw[15]), .A1(n44), .B0(enc_sboxw[15]), .B1(n47), 
        .Y(muxed_sboxw[15]) );
  INVX1 U23 ( .A(n75), .Y(n51) );
  INVX1 U24 ( .A(n69), .Y(n61) );
  INVX1 U25 ( .A(n71), .Y(n53) );
  INVX1 U26 ( .A(n70), .Y(n54) );
  INVX1 U27 ( .A(n70), .Y(n62) );
  INVX1 U28 ( .A(n64), .Y(n59) );
  INVX1 U29 ( .A(n67), .Y(n57) );
  INVX1 U30 ( .A(n72), .Y(n52) );
  INVX1 U31 ( .A(n63), .Y(n60) );
  INVX1 U32 ( .A(n66), .Y(n58) );
  INVX1 U33 ( .A(n69), .Y(n55) );
  INVX1 U34 ( .A(n68), .Y(n56) );
  INVX1 U35 ( .A(n47), .Y(n44) );
  INVX1 U36 ( .A(n46), .Y(n45) );
  BUFX2 U37 ( .A(n75), .Y(n73) );
  BUFX2 U38 ( .A(n78), .Y(n63) );
  BUFX2 U39 ( .A(n78), .Y(n64) );
  BUFX2 U40 ( .A(n76), .Y(n71) );
  BUFX2 U41 ( .A(n76), .Y(n70) );
  BUFX2 U42 ( .A(n77), .Y(n67) );
  BUFX2 U43 ( .A(n75), .Y(n72) );
  BUFX2 U44 ( .A(n77), .Y(n66) );
  BUFX2 U45 ( .A(n76), .Y(n69) );
  BUFX2 U46 ( .A(n78), .Y(n65) );
  BUFX2 U47 ( .A(n77), .Y(n68) );
  BUFX2 U48 ( .A(n64), .Y(n74) );
  BUFX2 U49 ( .A(n48), .Y(n46) );
  BUFX2 U50 ( .A(n49), .Y(n47) );
  BUFX2 U51 ( .A(n49), .Y(n48) );
  INVX1 U52 ( .A(n12), .Y(n81) );
  BUFX2 U53 ( .A(n79), .Y(n78) );
  BUFX2 U54 ( .A(n63), .Y(n75) );
  BUFX2 U55 ( .A(n64), .Y(n76) );
  BUFX2 U56 ( .A(n79), .Y(n77) );
  INVX1 U57 ( .A(n43), .Y(n49) );
  NOR2X1 U58 ( .A(n73), .B(n83), .Y(enc_next) );
  NAND2X1 U59 ( .A(n82), .B(n9), .Y(n12) );
  NOR2X1 U60 ( .A(n51), .B(n83), .Y(dec_next) );
  INVX1 U61 ( .A(n14), .Y(n82) );
  OAI211X1 U62 ( .A0(n11), .A1(n83), .B0(n13), .C0(n8), .Y(n14) );
  INVX1 U63 ( .A(n50), .Y(n79) );
  NAND2BX1 U64 ( .AN(n11), .B(init), .Y(n13) );
  AO22X1 U65 ( .A0(keymem_sboxw[10]), .A1(n44), .B0(enc_sboxw[10]), .B1(n47), 
        .Y(muxed_sboxw[10]) );
  AO22X1 U66 ( .A0(keymem_sboxw[14]), .A1(n44), .B0(enc_sboxw[14]), .B1(n47), 
        .Y(muxed_sboxw[14]) );
  AO22X1 U67 ( .A0(keymem_sboxw[13]), .A1(n44), .B0(enc_sboxw[13]), .B1(n47), 
        .Y(muxed_sboxw[13]) );
  BUFX2 U68 ( .A(n16), .Y(n43) );
  OAI21XL U69 ( .A0(aes_core_ctrl_reg[1]), .A1(n5), .B0(n13), .Y(n16) );
  NAND2X1 U70 ( .A(n5), .B(n4), .Y(n11) );
  AO22X1 U71 ( .A0(keymem_sboxw[0]), .A1(n44), .B0(enc_sboxw[0]), .B1(n46), 
        .Y(muxed_sboxw[0]) );
  AO22X1 U72 ( .A0(keymem_sboxw[2]), .A1(n16), .B0(enc_sboxw[2]), .B1(n48), 
        .Y(muxed_sboxw[2]) );
  AO22X1 U73 ( .A0(keymem_sboxw[5]), .A1(n43), .B0(enc_sboxw[5]), .B1(n48), 
        .Y(muxed_sboxw[5]) );
  AO22X1 U74 ( .A0(keymem_sboxw[4]), .A1(n43), .B0(enc_sboxw[4]), .B1(n48), 
        .Y(muxed_sboxw[4]) );
  AO22X1 U75 ( .A0(keymem_sboxw[1]), .A1(n45), .B0(n49), .B1(enc_sboxw[1]), 
        .Y(muxed_sboxw[1]) );
  AO22X1 U76 ( .A0(keymem_sboxw[3]), .A1(n43), .B0(enc_sboxw[3]), .B1(n48), 
        .Y(muxed_sboxw[3]) );
  AO22X1 U77 ( .A0(keymem_sboxw[6]), .A1(n16), .B0(enc_sboxw[6]), .B1(n48), 
        .Y(muxed_sboxw[6]) );
  AO22X1 U78 ( .A0(keymem_sboxw[7]), .A1(n16), .B0(enc_sboxw[7]), .B1(n46), 
        .Y(muxed_sboxw[7]) );
  AO22X1 U79 ( .A0(keymem_sboxw[20]), .A1(n45), .B0(enc_sboxw[20]), .B1(n46), 
        .Y(muxed_sboxw[20]) );
  AO22X1 U80 ( .A0(keymem_sboxw[19]), .A1(n45), .B0(enc_sboxw[19]), .B1(n46), 
        .Y(muxed_sboxw[19]) );
  AO22X1 U81 ( .A0(keymem_sboxw[21]), .A1(n45), .B0(enc_sboxw[21]), .B1(n46), 
        .Y(muxed_sboxw[21]) );
  AO22X1 U82 ( .A0(keymem_sboxw[29]), .A1(n16), .B0(enc_sboxw[29]), .B1(n48), 
        .Y(muxed_sboxw[29]) );
  AO22X1 U83 ( .A0(keymem_sboxw[28]), .A1(n16), .B0(enc_sboxw[28]), .B1(n48), 
        .Y(muxed_sboxw[28]) );
  AO22X1 U84 ( .A0(keymem_sboxw[27]), .A1(n45), .B0(enc_sboxw[27]), .B1(n49), 
        .Y(muxed_sboxw[27]) );
  AO22X1 U85 ( .A0(keymem_sboxw[26]), .A1(n45), .B0(enc_sboxw[26]), .B1(n49), 
        .Y(muxed_sboxw[26]) );
  AO22X1 U86 ( .A0(keymem_sboxw[18]), .A1(n44), .B0(enc_sboxw[18]), .B1(n47), 
        .Y(muxed_sboxw[18]) );
  AO22X1 U87 ( .A0(keymem_sboxw[24]), .A1(n45), .B0(enc_sboxw[24]), .B1(n46), 
        .Y(muxed_sboxw[24]) );
  AO22X1 U88 ( .A0(keymem_sboxw[25]), .A1(n45), .B0(enc_sboxw[25]), .B1(n46), 
        .Y(muxed_sboxw[25]) );
  AO22X1 U89 ( .A0(keymem_sboxw[16]), .A1(n44), .B0(enc_sboxw[16]), .B1(n47), 
        .Y(muxed_sboxw[16]) );
  AO22X1 U90 ( .A0(keymem_sboxw[17]), .A1(n44), .B0(enc_sboxw[17]), .B1(n47), 
        .Y(muxed_sboxw[17]) );
  AO22X1 U91 ( .A0(keymem_sboxw[30]), .A1(n16), .B0(enc_sboxw[30]), .B1(n46), 
        .Y(muxed_sboxw[30]) );
  AO22X1 U92 ( .A0(keymem_sboxw[22]), .A1(n45), .B0(enc_sboxw[22]), .B1(n49), 
        .Y(muxed_sboxw[22]) );
  AO22X1 U93 ( .A0(keymem_sboxw[23]), .A1(n45), .B0(enc_sboxw[23]), .B1(n49), 
        .Y(muxed_sboxw[23]) );
  AO22X1 U94 ( .A0(enc_round_nr[3]), .A1(n51), .B0(dec_round_nr[3]), .B1(n63), 
        .Y(muxed_round_nr[3]) );
  AO22X1 U95 ( .A0(enc_round_nr[1]), .A1(n51), .B0(dec_round_nr[1]), .B1(n67), 
        .Y(muxed_round_nr[1]) );
  AO22X1 U96 ( .A0(keymem_sboxw[31]), .A1(n16), .B0(enc_sboxw[31]), .B1(n46), 
        .Y(muxed_sboxw[31]) );
  AO22X1 U97 ( .A0(enc_round_nr[0]), .A1(n51), .B0(dec_round_nr[0]), .B1(n64), 
        .Y(muxed_round_nr[0]) );
  AO22X1 U98 ( .A0(enc_round_nr[2]), .A1(n51), .B0(dec_round_nr[2]), .B1(n66), 
        .Y(muxed_round_nr[2]) );
  NAND3X1 U99 ( .A(aes_core_ctrl_reg[0]), .B(n4), .C(key_ready), .Y(n9) );
  NAND3X1 U100 ( .A(n15), .B(n5), .C(aes_core_ctrl_reg[1]), .Y(n8) );
  AO22X1 U101 ( .A0(enc_ready), .A1(n51), .B0(dec_ready), .B1(n64), .Y(n15) );
  OAI21XL U102 ( .A0(n5), .A1(n12), .B0(n13), .Y(n20) );
  NAND3X1 U103 ( .A(n8), .B(n9), .C(n10), .Y(n18) );
  NAND2X1 U104 ( .A(ready), .B(n81), .Y(n10) );
  INVX1 U105 ( .A(next), .Y(n83) );
  OAI2BB1X1 U106 ( .A0N(result_valid), .A1N(n82), .B0(n8), .Y(n17) );
  OAI32X1 U107 ( .A0(n11), .A1(init), .A2(n81), .B0(n4), .B1(n12), .Y(n19) );
  AO22X1 U108 ( .A0(enc_new_block[7]), .A1(n61), .B0(dec_new_block[7]), .B1(
        n75), .Y(result[7]) );
  AO22X1 U109 ( .A0(enc_new_block[39]), .A1(n57), .B0(dec_new_block[39]), .B1(
        n67), .Y(result[39]) );
  AO22X1 U110 ( .A0(enc_new_block[15]), .A1(n55), .B0(dec_new_block[15]), .B1(
        n74), .Y(result[15]) );
  AO22X1 U111 ( .A0(enc_new_block[47]), .A1(n58), .B0(dec_new_block[47]), .B1(
        n65), .Y(result[47]) );
  AO22X1 U112 ( .A0(enc_new_block[6]), .A1(n60), .B0(dec_new_block[6]), .B1(
        n72), .Y(result[6]) );
  AO22X1 U113 ( .A0(enc_new_block[38]), .A1(n57), .B0(dec_new_block[38]), .B1(
        n66), .Y(result[38]) );
  AO22X1 U114 ( .A0(enc_new_block[14]), .A1(n54), .B0(dec_new_block[14]), .B1(
        n74), .Y(result[14]) );
  AO22X1 U115 ( .A0(enc_new_block[46]), .A1(n58), .B0(dec_new_block[46]), .B1(
        n65), .Y(result[46]) );
  AO22X1 U116 ( .A0(enc_new_block[5]), .A1(n50), .B0(dec_new_block[5]), .B1(
        n76), .Y(result[5]) );
  AO22X1 U117 ( .A0(enc_new_block[37]), .A1(n57), .B0(dec_new_block[37]), .B1(
        n68), .Y(result[37]) );
  AO22X1 U118 ( .A0(enc_new_block[13]), .A1(n54), .B0(dec_new_block[13]), .B1(
        n74), .Y(result[13]) );
  AO22X1 U119 ( .A0(enc_new_block[45]), .A1(n58), .B0(dec_new_block[45]), .B1(
        n72), .Y(result[45]) );
  AO22X1 U120 ( .A0(enc_new_block[4]), .A1(n58), .B0(dec_new_block[4]), .B1(
        n73), .Y(result[4]) );
  AO22X1 U121 ( .A0(enc_new_block[36]), .A1(n57), .B0(dec_new_block[36]), .B1(
        n65), .Y(result[36]) );
  AO22X1 U122 ( .A0(enc_new_block[12]), .A1(n54), .B0(dec_new_block[12]), .B1(
        n74), .Y(result[12]) );
  AO22X1 U123 ( .A0(enc_new_block[44]), .A1(n58), .B0(dec_new_block[44]), .B1(
        n71), .Y(result[44]) );
  AO22X1 U124 ( .A0(enc_new_block[3]), .A1(n57), .B0(dec_new_block[3]), .B1(
        n72), .Y(result[3]) );
  AO22X1 U125 ( .A0(enc_new_block[35]), .A1(n57), .B0(dec_new_block[35]), .B1(
        n68), .Y(result[35]) );
  AO22X1 U126 ( .A0(enc_new_block[11]), .A1(n53), .B0(dec_new_block[11]), .B1(
        n63), .Y(result[11]) );
  AO22X1 U127 ( .A0(enc_new_block[43]), .A1(n58), .B0(dec_new_block[43]), .B1(
        n70), .Y(result[43]) );
  AO22X1 U128 ( .A0(enc_new_block[2]), .A1(n56), .B0(dec_new_block[2]), .B1(
        n79), .Y(result[2]) );
  AO22X1 U129 ( .A0(enc_new_block[34]), .A1(n57), .B0(dec_new_block[34]), .B1(
        n79), .Y(result[34]) );
  AO22X1 U130 ( .A0(enc_new_block[10]), .A1(n52), .B0(dec_new_block[10]), .B1(
        n73), .Y(result[10]) );
  AO22X1 U131 ( .A0(enc_new_block[42]), .A1(n58), .B0(dec_new_block[42]), .B1(
        n71), .Y(result[42]) );
  AO22X1 U132 ( .A0(enc_new_block[0]), .A1(n51), .B0(dec_new_block[0]), .B1(
        n65), .Y(result[0]) );
  AO22X1 U133 ( .A0(enc_new_block[32]), .A1(n56), .B0(dec_new_block[32]), .B1(
        n79), .Y(result[32]) );
  AO22X1 U134 ( .A0(enc_new_block[8]), .A1(n62), .B0(dec_new_block[8]), .B1(
        n66), .Y(result[8]) );
  AO22X1 U135 ( .A0(enc_new_block[40]), .A1(n57), .B0(dec_new_block[40]), .B1(
        n70), .Y(result[40]) );
  AO22X1 U136 ( .A0(enc_new_block[1]), .A1(n55), .B0(dec_new_block[1]), .B1(
        n70), .Y(result[1]) );
  AO22X1 U137 ( .A0(enc_new_block[33]), .A1(n57), .B0(dec_new_block[33]), .B1(
        n68), .Y(result[33]) );
  AO22X1 U138 ( .A0(n50), .A1(enc_new_block[9]), .B0(dec_new_block[9]), .B1(
        n72), .Y(result[9]) );
  AO22X1 U139 ( .A0(enc_new_block[41]), .A1(n57), .B0(dec_new_block[41]), .B1(
        n69), .Y(result[41]) );
  AO22X1 U140 ( .A0(enc_new_block[71]), .A1(n60), .B0(dec_new_block[71]), .B1(
        n64), .Y(result[71]) );
  AO22X1 U141 ( .A0(enc_new_block[103]), .A1(n52), .B0(dec_new_block[103]), 
        .B1(n69), .Y(result[103]) );
  AO22X1 U142 ( .A0(enc_new_block[79]), .A1(n61), .B0(dec_new_block[79]), .B1(
        n69), .Y(result[79]) );
  AO22X1 U143 ( .A0(enc_new_block[111]), .A1(n52), .B0(dec_new_block[111]), 
        .B1(n73), .Y(result[111]) );
  AO22X1 U144 ( .A0(enc_new_block[70]), .A1(n60), .B0(dec_new_block[70]), .B1(
        n75), .Y(result[70]) );
  AO22X1 U145 ( .A0(enc_new_block[102]), .A1(n51), .B0(dec_new_block[102]), 
        .B1(n68), .Y(result[102]) );
  AO22X1 U146 ( .A0(enc_new_block[78]), .A1(n60), .B0(dec_new_block[78]), .B1(
        n71), .Y(result[78]) );
  AO22X1 U147 ( .A0(enc_new_block[110]), .A1(n52), .B0(dec_new_block[110]), 
        .B1(n73), .Y(result[110]) );
  AO22X1 U148 ( .A0(enc_new_block[69]), .A1(n59), .B0(dec_new_block[69]), .B1(
        n78), .Y(result[69]) );
  AO22X1 U149 ( .A0(enc_new_block[101]), .A1(n51), .B0(dec_new_block[101]), 
        .B1(n67), .Y(result[101]) );
  AO22X1 U150 ( .A0(enc_new_block[77]), .A1(n60), .B0(dec_new_block[77]), .B1(
        n70), .Y(result[77]) );
  AO22X1 U151 ( .A0(enc_new_block[109]), .A1(n52), .B0(dec_new_block[109]), 
        .B1(n73), .Y(result[109]) );
  AO22X1 U152 ( .A0(enc_new_block[68]), .A1(n59), .B0(dec_new_block[68]), .B1(
        n65), .Y(result[68]) );
  AO22X1 U153 ( .A0(enc_new_block[100]), .A1(n51), .B0(dec_new_block[100]), 
        .B1(n66), .Y(result[100]) );
  AO22X1 U154 ( .A0(enc_new_block[76]), .A1(n60), .B0(dec_new_block[76]), .B1(
        n69), .Y(result[76]) );
  AO22X1 U155 ( .A0(enc_new_block[108]), .A1(n52), .B0(dec_new_block[108]), 
        .B1(n73), .Y(result[108]) );
  AO22X1 U156 ( .A0(enc_new_block[67]), .A1(n59), .B0(dec_new_block[67]), .B1(
        n67), .Y(result[67]) );
  AO22X1 U157 ( .A0(enc_new_block[99]), .A1(n50), .B0(dec_new_block[99]), .B1(
        n71), .Y(result[99]) );
  AO22X1 U158 ( .A0(enc_new_block[75]), .A1(n60), .B0(dec_new_block[75]), .B1(
        n67), .Y(result[75]) );
  AO22X1 U159 ( .A0(enc_new_block[107]), .A1(n52), .B0(dec_new_block[107]), 
        .B1(n78), .Y(result[107]) );
  AO22X1 U160 ( .A0(enc_new_block[66]), .A1(n59), .B0(dec_new_block[66]), .B1(
        n77), .Y(result[66]) );
  AO22X1 U161 ( .A0(enc_new_block[98]), .A1(n50), .B0(dec_new_block[98]), .B1(
        n77), .Y(result[98]) );
  AO22X1 U162 ( .A0(enc_new_block[74]), .A1(n60), .B0(dec_new_block[74]), .B1(
        n66), .Y(result[74]) );
  AO22X1 U163 ( .A0(enc_new_block[106]), .A1(n52), .B0(dec_new_block[106]), 
        .B1(n72), .Y(result[106]) );
  AO22X1 U164 ( .A0(enc_new_block[64]), .A1(n59), .B0(dec_new_block[64]), .B1(
        n78), .Y(result[64]) );
  AO22X1 U165 ( .A0(enc_new_block[96]), .A1(n62), .B0(dec_new_block[96]), .B1(
        n73), .Y(result[96]) );
  AO22X1 U166 ( .A0(enc_new_block[72]), .A1(n60), .B0(dec_new_block[72]), .B1(
        n68), .Y(result[72]) );
  AO22X1 U167 ( .A0(enc_new_block[104]), .A1(n52), .B0(dec_new_block[104]), 
        .B1(n70), .Y(result[104]) );
  AO22X1 U168 ( .A0(enc_new_block[65]), .A1(n59), .B0(dec_new_block[65]), .B1(
        n75), .Y(result[65]) );
  AO22X1 U169 ( .A0(enc_new_block[97]), .A1(n50), .B0(dec_new_block[97]), .B1(
        n68), .Y(result[97]) );
  AO22X1 U170 ( .A0(enc_new_block[73]), .A1(n60), .B0(dec_new_block[73]), .B1(
        n79), .Y(result[73]) );
  AO22X1 U171 ( .A0(enc_new_block[105]), .A1(n52), .B0(dec_new_block[105]), 
        .B1(n71), .Y(result[105]) );
  BUFX2 U172 ( .A(encdec), .Y(n50) );
  AO22X1 U173 ( .A0(enc_new_block[87]), .A1(n61), .B0(dec_new_block[87]), .B1(
        n76), .Y(result[87]) );
  AO22X1 U174 ( .A0(enc_new_block[95]), .A1(n62), .B0(dec_new_block[95]), .B1(
        n72), .Y(result[95]) );
  AO22X1 U175 ( .A0(enc_new_block[86]), .A1(n61), .B0(dec_new_block[86]), .B1(
        n65), .Y(result[86]) );
  AO22X1 U176 ( .A0(enc_new_block[94]), .A1(n62), .B0(dec_new_block[94]), .B1(
        n71), .Y(result[94]) );
  AO22X1 U177 ( .A0(enc_new_block[85]), .A1(n61), .B0(dec_new_block[85]), .B1(
        n63), .Y(result[85]) );
  AO22X1 U178 ( .A0(enc_new_block[93]), .A1(n62), .B0(dec_new_block[93]), .B1(
        n79), .Y(result[93]) );
  AO22X1 U179 ( .A0(enc_new_block[84]), .A1(n61), .B0(dec_new_block[84]), .B1(
        n64), .Y(result[84]) );
  AO22X1 U180 ( .A0(enc_new_block[92]), .A1(n62), .B0(dec_new_block[92]), .B1(
        n78), .Y(result[92]) );
  AO22X1 U181 ( .A0(enc_new_block[83]), .A1(n61), .B0(dec_new_block[83]), .B1(
        n70), .Y(result[83]) );
  AO22X1 U182 ( .A0(enc_new_block[91]), .A1(n62), .B0(dec_new_block[91]), .B1(
        n75), .Y(result[91]) );
  AO22X1 U183 ( .A0(enc_new_block[82]), .A1(n61), .B0(dec_new_block[82]), .B1(
        n79), .Y(result[82]) );
  AO22X1 U184 ( .A0(enc_new_block[90]), .A1(n62), .B0(dec_new_block[90]), .B1(
        n76), .Y(result[90]) );
  AO22X1 U185 ( .A0(enc_new_block[80]), .A1(n61), .B0(dec_new_block[80]), .B1(
        n65), .Y(result[80]) );
  AO22X1 U186 ( .A0(enc_new_block[88]), .A1(n62), .B0(dec_new_block[88]), .B1(
        n69), .Y(result[88]) );
  AO22X1 U187 ( .A0(enc_new_block[81]), .A1(n61), .B0(dec_new_block[81]), .B1(
        n71), .Y(result[81]) );
  AO22X1 U188 ( .A0(enc_new_block[89]), .A1(n62), .B0(dec_new_block[89]), .B1(
        n77), .Y(result[89]) );
  AO22X1 U189 ( .A0(enc_new_block[119]), .A1(n53), .B0(dec_new_block[119]), 
        .B1(n64), .Y(result[119]) );
  AO22X1 U190 ( .A0(enc_new_block[127]), .A1(n54), .B0(dec_new_block[127]), 
        .B1(n74), .Y(result[127]) );
  AO22X1 U191 ( .A0(enc_new_block[118]), .A1(n53), .B0(dec_new_block[118]), 
        .B1(n66), .Y(result[118]) );
  AO22X1 U192 ( .A0(enc_new_block[126]), .A1(n54), .B0(dec_new_block[126]), 
        .B1(n74), .Y(result[126]) );
  AO22X1 U193 ( .A0(enc_new_block[117]), .A1(n53), .B0(dec_new_block[117]), 
        .B1(n68), .Y(result[117]) );
  AO22X1 U194 ( .A0(enc_new_block[125]), .A1(n54), .B0(dec_new_block[125]), 
        .B1(n74), .Y(result[125]) );
  AO22X1 U195 ( .A0(enc_new_block[116]), .A1(n53), .B0(dec_new_block[116]), 
        .B1(n79), .Y(result[116]) );
  AO22X1 U196 ( .A0(enc_new_block[124]), .A1(n54), .B0(dec_new_block[124]), 
        .B1(n74), .Y(result[124]) );
  AO22X1 U197 ( .A0(enc_new_block[115]), .A1(n53), .B0(dec_new_block[115]), 
        .B1(n78), .Y(result[115]) );
  AO22X1 U198 ( .A0(enc_new_block[123]), .A1(n54), .B0(dec_new_block[123]), 
        .B1(n74), .Y(result[123]) );
  AO22X1 U199 ( .A0(enc_new_block[114]), .A1(n53), .B0(dec_new_block[114]), 
        .B1(n75), .Y(result[114]) );
  AO22X1 U200 ( .A0(enc_new_block[122]), .A1(n54), .B0(dec_new_block[122]), 
        .B1(n74), .Y(result[122]) );
  AO22X1 U201 ( .A0(enc_new_block[120]), .A1(n53), .B0(dec_new_block[120]), 
        .B1(n76), .Y(result[120]) );
  AO22X1 U202 ( .A0(enc_new_block[113]), .A1(n53), .B0(dec_new_block[113]), 
        .B1(n63), .Y(result[113]) );
  AO22X1 U203 ( .A0(enc_new_block[121]), .A1(n54), .B0(dec_new_block[121]), 
        .B1(n77), .Y(result[121]) );
  AO22X1 U204 ( .A0(enc_new_block[112]), .A1(n53), .B0(dec_new_block[112]), 
        .B1(n73), .Y(result[112]) );
  AO22X1 U205 ( .A0(enc_new_block[23]), .A1(n55), .B0(dec_new_block[23]), .B1(
        n79), .Y(result[23]) );
  AO22X1 U206 ( .A0(enc_new_block[55]), .A1(n50), .B0(dec_new_block[55]), .B1(
        n66), .Y(result[55]) );
  AO22X1 U207 ( .A0(enc_new_block[22]), .A1(n55), .B0(dec_new_block[22]), .B1(
        n73), .Y(result[22]) );
  AO22X1 U208 ( .A0(enc_new_block[54]), .A1(n50), .B0(dec_new_block[54]), .B1(
        n65), .Y(result[54]) );
  AO22X1 U209 ( .A0(enc_new_block[21]), .A1(n55), .B0(dec_new_block[21]), .B1(
        n63), .Y(result[21]) );
  AO22X1 U210 ( .A0(enc_new_block[53]), .A1(n50), .B0(dec_new_block[53]), .B1(
        n71), .Y(result[53]) );
  AO22X1 U211 ( .A0(enc_new_block[20]), .A1(n55), .B0(dec_new_block[20]), .B1(
        n70), .Y(result[20]) );
  AO22X1 U212 ( .A0(enc_new_block[52]), .A1(n50), .B0(dec_new_block[52]), .B1(
        n63), .Y(result[52]) );
  AO22X1 U213 ( .A0(enc_new_block[19]), .A1(n55), .B0(dec_new_block[19]), .B1(
        n69), .Y(result[19]) );
  AO22X1 U214 ( .A0(enc_new_block[51]), .A1(encdec), .B0(dec_new_block[51]), 
        .B1(n69), .Y(result[51]) );
  AO22X1 U215 ( .A0(enc_new_block[18]), .A1(n55), .B0(dec_new_block[18]), .B1(
        n67), .Y(result[18]) );
  AO22X1 U216 ( .A0(enc_new_block[50]), .A1(n58), .B0(dec_new_block[50]), .B1(
        n67), .Y(result[50]) );
  AO22X1 U217 ( .A0(enc_new_block[16]), .A1(n55), .B0(dec_new_block[16]), .B1(
        n66), .Y(result[16]) );
  AO22X1 U218 ( .A0(enc_new_block[48]), .A1(n58), .B0(dec_new_block[48]), .B1(
        n66), .Y(result[48]) );
  AO22X1 U219 ( .A0(enc_new_block[17]), .A1(n55), .B0(dec_new_block[17]), .B1(
        n68), .Y(result[17]) );
  AO22X1 U220 ( .A0(enc_new_block[49]), .A1(n58), .B0(dec_new_block[49]), .B1(
        n68), .Y(result[49]) );
  AO22X1 U221 ( .A0(enc_new_block[31]), .A1(n56), .B0(dec_new_block[31]), .B1(
        n72), .Y(result[31]) );
  AO22X1 U222 ( .A0(enc_new_block[63]), .A1(n59), .B0(dec_new_block[63]), .B1(
        n76), .Y(result[63]) );
  AO22X1 U223 ( .A0(enc_new_block[30]), .A1(n56), .B0(dec_new_block[30]), .B1(
        n71), .Y(result[30]) );
  AO22X1 U224 ( .A0(enc_new_block[62]), .A1(n59), .B0(dec_new_block[62]), .B1(
        n67), .Y(result[62]) );
  AO22X1 U225 ( .A0(enc_new_block[29]), .A1(n56), .B0(dec_new_block[29]), .B1(
        n77), .Y(result[29]) );
  AO22X1 U226 ( .A0(enc_new_block[61]), .A1(n59), .B0(dec_new_block[61]), .B1(
        n65), .Y(result[61]) );
  AO22X1 U227 ( .A0(enc_new_block[28]), .A1(n56), .B0(dec_new_block[28]), .B1(
        n78), .Y(result[28]) );
  AO22X1 U228 ( .A0(enc_new_block[60]), .A1(n59), .B0(dec_new_block[60]), .B1(
        n77), .Y(result[60]) );
  AO22X1 U229 ( .A0(enc_new_block[27]), .A1(n56), .B0(dec_new_block[27]), .B1(
        n75), .Y(result[27]) );
  AO22X1 U230 ( .A0(enc_new_block[59]), .A1(encdec), .B0(dec_new_block[59]), 
        .B1(n67), .Y(result[59]) );
  AO22X1 U231 ( .A0(enc_new_block[26]), .A1(n56), .B0(dec_new_block[26]), .B1(
        n76), .Y(result[26]) );
  AO22X1 U232 ( .A0(enc_new_block[58]), .A1(encdec), .B0(dec_new_block[58]), 
        .B1(n63), .Y(result[58]) );
  AO22X1 U233 ( .A0(enc_new_block[24]), .A1(n56), .B0(dec_new_block[24]), .B1(
        n72), .Y(result[24]) );
  AO22X1 U234 ( .A0(enc_new_block[56]), .A1(encdec), .B0(dec_new_block[56]), 
        .B1(n64), .Y(result[56]) );
  AO22X1 U235 ( .A0(enc_new_block[25]), .A1(n56), .B0(dec_new_block[25]), .B1(
        n65), .Y(result[25]) );
  AO22X1 U236 ( .A0(enc_new_block[57]), .A1(encdec), .B0(dec_new_block[57]), 
        .B1(n72), .Y(result[57]) );
  INVX1 U237 ( .A(new_sboxw[15]), .Y(n2) );
  INVX1 U238 ( .A(new_sboxw[2]), .Y(n6) );
  INVX1 U239 ( .A(new_sboxw[3]), .Y(n21) );
  INVX1 U240 ( .A(new_sboxw[5]), .Y(n23) );
  INVX1 U241 ( .A(new_sboxw[13]), .Y(n25) );
  INVX1 U242 ( .A(new_sboxw[10]), .Y(n27) );
  INVX1 U243 ( .A(new_sboxw[7]), .Y(n29) );
  INVX1 U244 ( .A(new_sboxw[8]), .Y(n31) );
  INVX1 U245 ( .A(new_sboxw[4]), .Y(n33) );
  INVX1 U246 ( .A(new_sboxw[1]), .Y(n35) );
  INVX1 U247 ( .A(new_sboxw[14]), .Y(n37) );
  INVX1 U248 ( .A(new_sboxw[12]), .Y(n39) );
  INVX1 U249 ( .A(new_sboxw[9]), .Y(n41) );
endmodule


module display_DW01_inc_0 ( A, SUM );
  input [19:0] A;
  output [19:0] SUM;

  wire   [19:2] carry;

  ADDHXL U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[19]), .B(A[19]), .Y(SUM[19]) );
endmodule


module display ( clk, rst, data_in, sel, data_out );
  input [7:0] data_in;
  output [1:0] sel;
  output [6:0] data_out;
  input clk, rst;
  wire   N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19,
         N20, N21, N22, N23, N24, clkout, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47,
         scan_cnt, n78, n14, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n61, n62, n65, n1, n2, n3, n4, n5, n6, n8, n9, n10, n11,
         n12, n13, n15, n16, n17, n18, n59, n60, n63, n64, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77;
  wire   [19:0] cnt;
  assign sel[1] = scan_cnt;

  display_DW01_inc_0 add_29 ( .A(cnt), .SUM({N24, N23, N22, N21, N20, N19, N18, 
        N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5}) );
  DFFQX1 clkout_reg ( .D(n65), .CK(clk), .Q(clkout) );
  DFFRX1 \cnt_reg[18]  ( .D(N46), .CK(clk), .RN(rst), .Q(cnt[18]) );
  DFFRX1 \cnt_reg[16]  ( .D(N44), .CK(clk), .RN(rst), .Q(cnt[16]) );
  DFFRX1 \cnt_reg[19]  ( .D(N47), .CK(clk), .RN(n15), .Q(cnt[19]), .QN(n3) );
  DFFRX1 \cnt_reg[17]  ( .D(N45), .CK(clk), .RN(rst), .Q(cnt[17]) );
  DFFRX1 \cnt_reg[14]  ( .D(N42), .CK(clk), .RN(n15), .Q(cnt[14]) );
  DFFRX1 \cnt_reg[15]  ( .D(N43), .CK(clk), .RN(n15), .Q(cnt[15]), .QN(n2) );
  DFFRX1 \cnt_reg[12]  ( .D(N40), .CK(clk), .RN(n15), .Q(cnt[12]), .QN(n5) );
  DFFRX1 \cnt_reg[13]  ( .D(N41), .CK(clk), .RN(n15), .Q(cnt[13]), .QN(n1) );
  DFFRX1 \cnt_reg[6]  ( .D(N34), .CK(clk), .RN(n13), .Q(cnt[6]) );
  DFFRX1 \cnt_reg[11]  ( .D(N39), .CK(clk), .RN(n15), .Q(cnt[11]), .QN(n10) );
  DFFRX1 \cnt_reg[5]  ( .D(N33), .CK(clk), .RN(n13), .Q(cnt[5]) );
  DFFRX1 \cnt_reg[8]  ( .D(N36), .CK(clk), .RN(n13), .Q(cnt[8]) );
  DFFRX1 \cnt_reg[7]  ( .D(N35), .CK(clk), .RN(n13), .Q(cnt[7]) );
  DFFRX1 \cnt_reg[9]  ( .D(N37), .CK(clk), .RN(n13), .Q(cnt[9]) );
  DFFRX1 \cnt_reg[10]  ( .D(N38), .CK(clk), .RN(n15), .Q(cnt[10]), .QN(n4) );
  DFFRX1 \cnt_reg[3]  ( .D(N31), .CK(clk), .RN(n13), .Q(cnt[3]) );
  DFFRX1 \cnt_reg[1]  ( .D(N29), .CK(clk), .RN(n13), .Q(cnt[1]) );
  DFFRX1 \cnt_reg[4]  ( .D(N32), .CK(clk), .RN(n13), .Q(cnt[4]) );
  DFFRX1 \cnt_reg[2]  ( .D(N30), .CK(clk), .RN(n13), .Q(cnt[2]) );
  DFFRX1 \cnt_reg[0]  ( .D(N28), .CK(clk), .RN(n15), .Q(cnt[0]), .QN(n11) );
  DFFRX1 scan_cnt_reg ( .D(sel[0]), .CK(clkout), .RN(n15), .Q(scan_cnt), .QN(
        n78) );
  OAI221X1 U3 ( .A0(scan_cnt), .A1(n53), .B0(sel[0]), .B1(n54), .C0(n35), .Y(
        data_out[0]) );
  OAI221X1 U4 ( .A0(scan_cnt), .A1(n47), .B0(sel[0]), .B1(n48), .C0(n35), .Y(
        data_out[1]) );
  OAI221X1 U5 ( .A0(scan_cnt), .A1(n43), .B0(sel[0]), .B1(n44), .C0(n28), .Y(
        data_out[2]) );
  OAI221X1 U6 ( .A0(scan_cnt), .A1(n33), .B0(sel[0]), .B1(n34), .C0(n35), .Y(
        data_out[4]) );
  INVXL U7 ( .A(n78), .Y(n6) );
  INVX16 U8 ( .A(n6), .Y(sel[0]) );
  NOR2X1 U9 ( .A(data_in[0]), .B(scan_cnt), .Y(n26) );
  BUFX2 U10 ( .A(rst), .Y(n13) );
  BUFX2 U11 ( .A(rst), .Y(n15) );
  NOR2X1 U12 ( .A(n76), .B(data_in[1]), .Y(n42) );
  INVX1 U13 ( .A(data_in[1]), .Y(n71) );
  NOR2X1 U14 ( .A(n77), .B(data_in[1]), .Y(n32) );
  OAI2BB2XL U15 ( .B0(data_in[0]), .B1(n76), .A0N(n77), .A1N(n42), .Y(n57) );
  OR2X1 U16 ( .A(data_in[0]), .B(n71), .Y(n46) );
  INVX1 U17 ( .A(n12), .Y(n63) );
  OAI211X1 U18 ( .A0(n38), .A1(n70), .B0(n19), .C0(n39), .Y(data_out[3]) );
  INVX1 U19 ( .A(n26), .Y(n70) );
  AOI221XL U20 ( .A0(n77), .A1(n76), .B0(data_in[2]), .B1(data_in[1]), .C0(n42), .Y(n38) );
  INVX1 U21 ( .A(data_in[5]), .Y(n74) );
  NAND2X1 U22 ( .A(data_in[7]), .B(n74), .Y(n41) );
  AOI222XL U23 ( .A0(n24), .A1(data_in[0]), .B0(n25), .B1(data_in[4]), .C0(n22), .C1(n40), .Y(n39) );
  OAI221XL U24 ( .A0(n74), .A1(n73), .B0(data_in[7]), .B1(data_in[6]), .C0(n41), .Y(n40) );
  NAND2X1 U25 ( .A(data_in[2]), .B(n52), .Y(n51) );
  XOR2X1 U26 ( .A(data_in[1]), .B(data_in[0]), .Y(n52) );
  NAND3X1 U27 ( .A(n28), .B(n69), .C(n29), .Y(data_out[5]) );
  AOI22X1 U28 ( .A0(n74), .A1(n22), .B0(n26), .B1(n71), .Y(n29) );
  OAI22XL U29 ( .A0(data_in[4]), .A1(n72), .B0(data_in[6]), .B1(n41), .Y(n55)
         );
  NAND4X1 U30 ( .A(n19), .B(n20), .C(n69), .D(n21), .Y(data_out[6]) );
  NAND2X1 U31 ( .A(n26), .B(n27), .Y(n20) );
  AOI211X1 U32 ( .A0(n22), .A1(n23), .B0(n24), .C0(n25), .Y(n21) );
  AOI22X1 U33 ( .A0(n73), .A1(n22), .B0(n77), .B1(n26), .Y(n35) );
  NOR2X1 U34 ( .A(n77), .B(data_in[3]), .Y(n27) );
  NAND2X1 U35 ( .A(data_in[6]), .B(n50), .Y(n49) );
  XOR2X1 U36 ( .A(data_in[5]), .B(data_in[4]), .Y(n50) );
  INVX1 U37 ( .A(data_in[6]), .Y(n73) );
  INVX1 U38 ( .A(data_in[2]), .Y(n77) );
  NOR2X1 U39 ( .A(data_in[5]), .B(data_in[6]), .Y(n36) );
  NOR2X1 U40 ( .A(data_in[1]), .B(data_in[2]), .Y(n37) );
  NOR2X1 U41 ( .A(n73), .B(data_in[7]), .Y(n23) );
  NOR2X1 U42 ( .A(n73), .B(data_in[5]), .Y(n31) );
  INVX1 U43 ( .A(data_in[3]), .Y(n76) );
  NAND2X1 U44 ( .A(n75), .B(data_in[5]), .Y(n45) );
  INVX1 U45 ( .A(data_in[7]), .Y(n72) );
  AOI2BB1X1 U46 ( .A0N(n72), .A1N(data_in[6]), .B0(n74), .Y(n56) );
  AOI2BB1X1 U47 ( .A0N(n76), .A1N(data_in[2]), .B0(n71), .Y(n58) );
  INVX1 U48 ( .A(data_in[4]), .Y(n75) );
  NOR2BX1 U49 ( .AN(N21), .B(n63), .Y(N44) );
  NOR2BX1 U50 ( .AN(N23), .B(n63), .Y(N46) );
  AND2X2 U51 ( .A(N22), .B(n12), .Y(N45) );
  NOR2BX1 U52 ( .AN(N18), .B(n63), .Y(N41) );
  NOR2BX1 U53 ( .AN(N15), .B(n63), .Y(N38) );
  NOR2BX1 U54 ( .AN(N17), .B(n63), .Y(N40) );
  NOR2BX1 U55 ( .AN(N20), .B(n63), .Y(N43) );
  BUFX2 U56 ( .A(n14), .Y(n12) );
  AND2X2 U57 ( .A(N19), .B(n12), .Y(N42) );
  AND2X2 U58 ( .A(N14), .B(n12), .Y(N37) );
  AND2X2 U59 ( .A(N16), .B(n12), .Y(N39) );
  NOR2BX1 U60 ( .AN(N10), .B(n63), .Y(N33) );
  AND2X2 U61 ( .A(N7), .B(n12), .Y(N30) );
  AND2X2 U62 ( .A(N9), .B(n14), .Y(N32) );
  AND2X2 U63 ( .A(N6), .B(n12), .Y(N29) );
  AND2X2 U64 ( .A(N8), .B(n14), .Y(N31) );
  AND2X2 U65 ( .A(N12), .B(n14), .Y(N35) );
  AND2X2 U66 ( .A(N13), .B(n14), .Y(N36) );
  AND2X2 U67 ( .A(N11), .B(n14), .Y(N34) );
  AOI22XL U68 ( .A0(sel[0]), .A1(n27), .B0(scan_cnt), .B1(n23), .Y(n28) );
  NOR2XL U69 ( .A(sel[0]), .B(data_in[4]), .Y(n22) );
  NOR3XL U70 ( .A(sel[0]), .B(data_in[6]), .C(n74), .Y(n25) );
  AOI211X1 U71 ( .A0(n23), .A1(data_in[4]), .B0(n55), .C0(n56), .Y(n54) );
  AOI211X1 U72 ( .A0(n27), .A1(data_in[0]), .B0(n57), .C0(n58), .Y(n53) );
  AOI2BB2X1 U73 ( .B0(n49), .B1(n72), .A0N(n41), .A1N(n75), .Y(n48) );
  AOI22X1 U74 ( .A0(n42), .A1(data_in[0]), .B0(n51), .B1(n76), .Y(n47) );
  AOI222XL U75 ( .A0(data_in[7]), .A1(n73), .B0(n45), .B1(n72), .C0(data_in[4]), .C1(n74), .Y(n44) );
  AOI222XL U76 ( .A0(data_in[3]), .A1(n77), .B0(n46), .B1(n76), .C0(data_in[0]), .C1(n71), .Y(n43) );
  OA22X1 U77 ( .A0(n74), .A1(data_in[4]), .B0(n36), .B1(n72), .Y(n34) );
  OA22X1 U78 ( .A0(n71), .A1(data_in[0]), .B0(n37), .B1(n76), .Y(n33) );
  INVX1 U79 ( .A(n30), .Y(n69) );
  OAI33XL U80 ( .A0(n72), .A1(sel[0]), .A2(n31), .B0(n76), .B1(scan_cnt), .B2(
        n32), .Y(n30) );
  NOR3X1 U81 ( .A(data_in[2]), .B(scan_cnt), .C(n71), .Y(n24) );
  AOI33XL U82 ( .A0(data_in[4]), .A1(scan_cnt), .A2(n31), .B0(data_in[0]), 
        .B1(sel[0]), .B2(n32), .Y(n19) );
  NAND4BX1 U83 ( .AN(n59), .B(n61), .C(n3), .D(n13), .Y(n68) );
  NAND3BX1 U84 ( .AN(cnt[16]), .B(n1), .C(n4), .Y(n59) );
  NOR2BX1 U85 ( .AN(N24), .B(n63), .Y(N47) );
  OAI31XL U86 ( .A0(n68), .A1(n67), .A2(n66), .B0(n64), .Y(n65) );
  NAND3BX1 U87 ( .AN(n5), .B(cnt[5]), .C(cnt[15]), .Y(n66) );
  NAND3BX1 U88 ( .AN(n8), .B(cnt[18]), .C(n62), .Y(n67) );
  AO21X1 U89 ( .A0(n15), .A1(n63), .B0(n60), .Y(n64) );
  OR4X1 U90 ( .A(cnt[5]), .B(cnt[12]), .C(n18), .D(n17), .Y(n14) );
  NAND3BX1 U91 ( .AN(cnt[18]), .B(n61), .C(n2), .Y(n18) );
  NAND4BX1 U92 ( .AN(n16), .B(cnt[10]), .C(cnt[16]), .D(cnt[13]), .Y(n17) );
  NAND3BX1 U93 ( .AN(n8), .B(cnt[19]), .C(n62), .Y(n16) );
  NAND4X1 U94 ( .A(cnt[6]), .B(n9), .C(n10), .D(n11), .Y(n8) );
  AND3X2 U95 ( .A(cnt[8]), .B(cnt[7]), .C(cnt[9]), .Y(n9) );
  NOR3X1 U96 ( .A(cnt[14]), .B(cnt[1]), .C(cnt[17]), .Y(n61) );
  NOR3X1 U97 ( .A(cnt[2]), .B(cnt[4]), .C(cnt[3]), .Y(n62) );
  AND2X2 U98 ( .A(N5), .B(n12), .Y(N28) );
  INVX1 U99 ( .A(clkout), .Y(n60) );
endmodule


module aes ( XIN, XOUT, CLK, RST, DATA_7, DATA_6, DATA_5, DATA_4, DATA_3, 
        DATA_2, DATA_1, DATA_0, POS_1, POS_0, SEG_6, SEG_5, SEG_4, SEG_3, 
        SEG_2, SEG_1, SEG_0, FLAG, ENC_DEC, KEY_LEN, PHASE_2, PHASE_1, PHASE_0
 );
  input XIN, CLK, RST;
  output XOUT, POS_1, POS_0, SEG_6, SEG_5, SEG_4, SEG_3, SEG_2, SEG_1, SEG_0,
         FLAG, ENC_DEC, KEY_LEN, PHASE_2, PHASE_1, PHASE_0;
  inout DATA_7,  DATA_6,  DATA_5,  DATA_4,  DATA_3,  DATA_2,  DATA_1,  DATA_0;
  wire   sysclock, clock, reset, _8_net_, ready, result_valid, encdec, keylen,
         init, next, N57, N58, N94, N97, N98, N99, N100, N108, n8, n9, n10,
         n11, n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n121, n123, n124, n125, n127, n128, n129, n130, n131,
         n132, n133, n137, n138, n140, n142, n143, n145, n146, n147, n148,
         n150, n151, n152, n153, n154, n155, n157, n159, n160, n162, n164,
         n165, n167, n168, n170, n171, n172, n174, n175, n177, n178, n180,
         n181, n183, n185, n186, n188, n190, n192, n194, n196, n198, n200,
         n202, n204, n205, n207, n209, n211, n213, n214, n216, n218, n220,
         n222, n223, n224, n226, n227, n232, n233, n235, n236, n237, n238,
         n239, n241, n244, n249, n255, n256, n258, n260, n263, n266, n267,
         n269, n270, n272, n274, n276, n277, n279, n280, n282, n284, n285,
         n288, n291, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, \r80/carry[4] , \r80/carry[3] , \r80/carry[2] ,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332;
  wire   [7:0] result_reg;
  wire   [7:0] data;
  wire   [1:0] pos;
  wire   [6:0] seg;
  wire   [2:0] phase;
  wire   [7:0] display_data;
  wire   [255:0] key;
  wire   [127:0] block;
  wire   [127:0] result;
  wire   [2:0] next_status;
  wire   [4:0] cnt_32;
  tri   DATA_7;
  tri   DATA_6;
  tri   DATA_5;
  tri   DATA_4;
  tri   DATA_3;
  tri   DATA_2;
  tri   DATA_1;
  tri   DATA_0;

  PX3W SCLK_PAD ( .XIN(XIN), .XOUT(XOUT), .XC(sysclock) );
  PIDW CLK_PAD ( .PAD(CLK), .C(clock) );
  PIUW RST_PAD ( .PAD(RST), .C(reset) );
  PBD20W DATA_7_PAD ( .I(result_reg[7]), .OEN(n1191), .PAD(DATA_7), .C(data[7]) );
  PBD20W DATA_6_PAD ( .I(result_reg[6]), .OEN(n1191), .PAD(DATA_6), .C(data[6]) );
  PBD20W DATA_5_PAD ( .I(result_reg[5]), .OEN(n1190), .PAD(DATA_5), .C(data[5]) );
  PBD20W DATA_4_PAD ( .I(result_reg[4]), .OEN(n1190), .PAD(DATA_4), .C(data[4]) );
  PBD20W DATA_3_PAD ( .I(result_reg[3]), .OEN(n1189), .PAD(DATA_3), .C(data[3]) );
  PBD20W DATA_2_PAD ( .I(result_reg[2]), .OEN(n1189), .PAD(DATA_2), .C(data[2]) );
  PBD20W DATA_1_PAD ( .I(result_reg[1]), .OEN(n1189), .PAD(DATA_1), .C(data[1]) );
  PBD20W DATA_0_PAD ( .I(result_reg[0]), .OEN(n1190), .PAD(DATA_0), .C(data[0]) );
  PO20W POS_1_PAD ( .I(pos[1]), .PAD(POS_1) );
  PO20W POS_0_PAD ( .I(pos[0]), .PAD(POS_0) );
  PO20W SEG_6_PAD ( .I(seg[6]), .PAD(SEG_6) );
  PO20W SEG_5_PAD ( .I(seg[5]), .PAD(SEG_5) );
  PO20W SEG_4_PAD ( .I(seg[4]), .PAD(SEG_4) );
  PO20W SEG_3_PAD ( .I(seg[3]), .PAD(SEG_3) );
  PO20W SEG_2_PAD ( .I(seg[2]), .PAD(SEG_2) );
  PO20W SEG_1_PAD ( .I(seg[1]), .PAD(SEG_1) );
  PO20W SEG_0_PAD ( .I(seg[0]), .PAD(SEG_0) );
  PO20W FLAG_PAD ( .I(_8_net_), .PAD(FLAG) );
  PO20W ENC_DEC_PAD ( .I(encdec), .PAD(ENC_DEC) );
  PO20W KEY_LEN_PAD ( .I(keylen), .PAD(KEY_LEN) );
  PO20W PHASE_2_PAD ( .I(phase[2]), .PAD(PHASE_2) );
  PO20W PHASE_1_PAD ( .I(phase[1]), .PAD(PHASE_1) );
  PO20W PHASE_0_PAD ( .I(phase[0]), .PAD(PHASE_0) );
  aes_core aes_core ( .clk(sysclock), .reset_n(reset), .encdec(encdec), .init(
        init), .next(next), .ready(ready), .key(key), .keylen(n1102), .block(
        block), .result(result), .result_valid(result_valid) );
  display display ( .clk(sysclock), .rst(n1268), .data_in(display_data), .sel(
        pos), .data_out(seg) );
  DFFRX1 \key_reg[54]  ( .D(n747), .CK(n1304), .RN(n1270), .Q(key[54]), .QN(
        n355) );
  DFFRX1 \key_reg[78]  ( .D(n755), .CK(n1307), .RN(n1264), .Q(key[78]), .QN(
        n363) );
  DFFRX1 drive_reg ( .D(n1080), .CK(n1273), .RN(n1259), .Q(n1090), .QN(n1089)
         );
  DFFRX1 \block_reg[0]  ( .D(n1088), .CK(n1273), .RN(n1259), .Q(block[0]), 
        .QN(n685) );
  DFFRX1 \block_reg[41]  ( .D(n1072), .CK(n1274), .RN(n1260), .Q(block[41]), 
        .QN(n674) );
  DFFRX1 \block_reg[105]  ( .D(n1071), .CK(n1274), .RN(n1267), .Q(block[105]), 
        .QN(n673) );
  DFFRX1 \block_reg[9]  ( .D(n1054), .CK(n1276), .RN(n1272), .Q(block[9]), 
        .QN(n656) );
  DFFRX1 \block_reg[73]  ( .D(n1053), .CK(n1276), .RN(n1271), .Q(block[73]), 
        .QN(n655) );
  DFFRX1 \block_reg[33]  ( .D(n1048), .CK(n1277), .RN(n1262), .Q(block[33]), 
        .QN(n650) );
  DFFRX1 \block_reg[97]  ( .D(n1047), .CK(n1277), .RN(n1271), .Q(block[97]), 
        .QN(n649) );
  DFFRX1 \block_reg[49]  ( .D(n1042), .CK(n1277), .RN(n1261), .Q(block[49]), 
        .QN(n644) );
  DFFRX1 \block_reg[113]  ( .D(n1041), .CK(n1277), .RN(n1264), .Q(block[113]), 
        .QN(n643) );
  DFFRX1 \block_reg[17]  ( .D(n1036), .CK(n1278), .RN(n1228), .Q(block[17]), 
        .QN(n638) );
  DFFRX1 \block_reg[81]  ( .D(n1035), .CK(n1278), .RN(n1228), .Q(block[81]), 
        .QN(n637) );
  DFFRX1 \block_reg[1]  ( .D(n1030), .CK(n1278), .RN(n1229), .Q(block[1]), 
        .QN(n632) );
  DFFRX1 \block_reg[65]  ( .D(n1029), .CK(n1278), .RN(n1229), .Q(block[65]), 
        .QN(n631) );
  DFFRX1 \block_reg[104]  ( .D(n1026), .CK(n1279), .RN(n1229), .Q(block[104]), 
        .QN(n629) );
  DFFRX1 \block_reg[72]  ( .D(n1024), .CK(n1279), .RN(n1229), .Q(block[72]), 
        .QN(n627) );
  DFFRX1 \block_reg[40]  ( .D(n1022), .CK(n1279), .RN(n1229), .Q(block[40]), 
        .QN(n625) );
  DFFRX1 \block_reg[8]  ( .D(n1020), .CK(n1279), .RN(n1230), .Q(block[8]), 
        .QN(n623) );
  DFFRX1 \block_reg[16]  ( .D(n1019), .CK(n1279), .RN(n1230), .Q(block[16]), 
        .QN(n622) );
  DFFRX1 \block_reg[32]  ( .D(n1018), .CK(n1280), .RN(n1230), .Q(block[32]), 
        .QN(n621) );
  DFFRX1 \block_reg[48]  ( .D(n1017), .CK(n1280), .RN(n1230), .Q(block[48]), 
        .QN(n620) );
  DFFRX1 \block_reg[64]  ( .D(n1016), .CK(n1280), .RN(n1230), .Q(block[64]), 
        .QN(n619) );
  DFFRX1 \block_reg[80]  ( .D(n1015), .CK(n1280), .RN(n1230), .Q(block[80]), 
        .QN(n618) );
  DFFRX1 \block_reg[96]  ( .D(n1014), .CK(n1280), .RN(n1230), .Q(block[96]), 
        .QN(n617) );
  DFFRX1 \block_reg[112]  ( .D(n1013), .CK(n1280), .RN(n1230), .Q(block[112]), 
        .QN(n616) );
  DFFRX1 \block_reg[106]  ( .D(n977), .CK(n1284), .RN(n1234), .Q(block[106]), 
        .QN(n581) );
  DFFRX1 \block_reg[74]  ( .D(n975), .CK(n1284), .RN(n1234), .Q(block[74]), 
        .QN(n579) );
  DFFRX1 \block_reg[42]  ( .D(n973), .CK(n1284), .RN(n1234), .Q(block[42]), 
        .QN(n577) );
  DFFRX1 \block_reg[10]  ( .D(n971), .CK(n1284), .RN(n1234), .Q(block[10]), 
        .QN(n575) );
  DFFRX1 \block_reg[2]  ( .D(n970), .CK(n1284), .RN(n1235), .Q(block[2]), .QN(
        n574) );
  DFFRX1 \block_reg[18]  ( .D(n969), .CK(n1284), .RN(n1235), .Q(block[18]), 
        .QN(n573) );
  DFFRX1 \block_reg[34]  ( .D(n968), .CK(n1285), .RN(n1235), .Q(block[34]), 
        .QN(n572) );
  DFFRX1 \block_reg[50]  ( .D(n967), .CK(n1285), .RN(n1235), .Q(block[50]), 
        .QN(n571) );
  DFFRX1 \block_reg[66]  ( .D(n966), .CK(n1285), .RN(n1235), .Q(block[66]), 
        .QN(n570) );
  DFFRX1 \block_reg[82]  ( .D(n965), .CK(n1285), .RN(n1235), .Q(block[82]), 
        .QN(n569) );
  DFFRX1 \block_reg[98]  ( .D(n964), .CK(n1285), .RN(n1235), .Q(block[98]), 
        .QN(n568) );
  DFFRX1 \block_reg[114]  ( .D(n963), .CK(n1285), .RN(n1235), .Q(block[114]), 
        .QN(n567) );
  DFFRX1 \block_reg[107]  ( .D(n928), .CK(n1289), .RN(n1239), .Q(block[107]), 
        .QN(n533) );
  DFFRX1 \block_reg[75]  ( .D(n926), .CK(n1289), .RN(n1239), .Q(block[75]), 
        .QN(n531) );
  DFFRX1 \block_reg[43]  ( .D(n924), .CK(n1289), .RN(n1239), .Q(block[43]), 
        .QN(n529) );
  DFFRX1 \block_reg[11]  ( .D(n922), .CK(n1289), .RN(n1239), .Q(block[11]), 
        .QN(n527) );
  DFFRX1 \block_reg[3]  ( .D(n921), .CK(n1289), .RN(n1239), .Q(block[3]), .QN(
        n526) );
  DFFRX1 \block_reg[19]  ( .D(n920), .CK(n1289), .RN(n1240), .Q(block[19]), 
        .QN(n525) );
  DFFRX1 \block_reg[35]  ( .D(n919), .CK(n1289), .RN(n1240), .Q(block[35]), 
        .QN(n524) );
  DFFRX1 \block_reg[51]  ( .D(n918), .CK(n1290), .RN(n1240), .Q(block[51]), 
        .QN(n523) );
  DFFRX1 \block_reg[67]  ( .D(n917), .CK(n1290), .RN(n1240), .Q(block[67]), 
        .QN(n522) );
  DFFRX1 \block_reg[83]  ( .D(n916), .CK(n1290), .RN(n1240), .Q(block[83]), 
        .QN(n521) );
  DFFRX1 \block_reg[99]  ( .D(n915), .CK(n1290), .RN(n1240), .Q(block[99]), 
        .QN(n520) );
  DFFRX1 \block_reg[115]  ( .D(n914), .CK(n1290), .RN(n1240), .Q(block[115]), 
        .QN(n519) );
  DFFRX1 \block_reg[108]  ( .D(n879), .CK(n1293), .RN(n1244), .Q(block[108]), 
        .QN(n485) );
  DFFRX1 \block_reg[76]  ( .D(n877), .CK(n1294), .RN(n1244), .Q(block[76]), 
        .QN(n483) );
  DFFRX1 \block_reg[44]  ( .D(n875), .CK(n1294), .RN(n1244), .Q(block[44]), 
        .QN(n481) );
  DFFRX1 \block_reg[12]  ( .D(n873), .CK(n1294), .RN(n1244), .Q(block[12]), 
        .QN(n479) );
  DFFRX1 \block_reg[4]  ( .D(n872), .CK(n1294), .RN(n1244), .Q(block[4]), .QN(
        n478) );
  DFFRX1 \block_reg[20]  ( .D(n871), .CK(n1294), .RN(n1244), .Q(block[20]), 
        .QN(n477) );
  DFFRX1 \block_reg[36]  ( .D(n870), .CK(n1294), .RN(n1245), .Q(block[36]), 
        .QN(n476) );
  DFFRX1 \block_reg[52]  ( .D(n869), .CK(n1294), .RN(n1245), .Q(block[52]), 
        .QN(n475) );
  DFFRX1 \block_reg[68]  ( .D(n868), .CK(n1295), .RN(n1245), .Q(block[68]), 
        .QN(n474) );
  DFFRX1 \block_reg[84]  ( .D(n867), .CK(n1295), .RN(n1245), .Q(block[84]), 
        .QN(n473) );
  DFFRX1 \block_reg[100]  ( .D(n866), .CK(n1295), .RN(n1245), .Q(block[100]), 
        .QN(n472) );
  DFFRX1 \block_reg[116]  ( .D(n865), .CK(n1295), .RN(n1245), .Q(block[116]), 
        .QN(n471) );
  DFFRX1 \block_reg[109]  ( .D(n830), .CK(n1298), .RN(reset), .Q(block[109]), 
        .QN(n437) );
  DFFRX1 \block_reg[77]  ( .D(n828), .CK(n1299), .RN(reset), .Q(block[77]), 
        .QN(n435) );
  DFFRX1 \block_reg[45]  ( .D(n826), .CK(n1299), .RN(reset), .Q(block[45]), 
        .QN(n433) );
  DFFRX1 \block_reg[13]  ( .D(n824), .CK(n1299), .RN(n1271), .Q(block[13]), 
        .QN(n431) );
  DFFRX1 \block_reg[5]  ( .D(n823), .CK(n1299), .RN(n1261), .Q(block[5]), .QN(
        n430) );
  DFFRX1 \block_reg[21]  ( .D(n822), .CK(n1299), .RN(n1269), .Q(block[21]), 
        .QN(n429) );
  DFFRX1 \block_reg[37]  ( .D(n821), .CK(n1299), .RN(n1259), .Q(block[37]), 
        .QN(n428) );
  DFFRX1 \block_reg[53]  ( .D(n820), .CK(n1299), .RN(n1248), .Q(block[53]), 
        .QN(n427) );
  DFFRX1 \block_reg[69]  ( .D(n819), .CK(n1299), .RN(n1248), .Q(block[69]), 
        .QN(n426) );
  DFFRX1 \block_reg[85]  ( .D(n818), .CK(n1300), .RN(n1248), .Q(block[85]), 
        .QN(n425) );
  DFFRX1 \block_reg[101]  ( .D(n817), .CK(n1300), .RN(n1248), .Q(block[101]), 
        .QN(n424) );
  DFFRX1 \block_reg[117]  ( .D(n816), .CK(n1300), .RN(n1248), .Q(block[117]), 
        .QN(n423) );
  DFFRX1 \block_reg[110]  ( .D(n781), .CK(n1311), .RN(n1251), .Q(block[110]), 
        .QN(n389) );
  DFFRX1 \block_reg[78]  ( .D(n779), .CK(n1310), .RN(n1252), .Q(block[78]), 
        .QN(n387) );
  DFFRX1 \block_reg[46]  ( .D(n777), .CK(n1306), .RN(n1252), .Q(block[46]), 
        .QN(n385) );
  DFFRX1 \block_reg[14]  ( .D(n775), .CK(clock), .RN(n1252), .Q(block[14]), 
        .QN(n383) );
  DFFRX1 \block_reg[6]  ( .D(n774), .CK(clock), .RN(n1252), .Q(block[6]), .QN(
        n382) );
  DFFRX1 \block_reg[22]  ( .D(n773), .CK(n1312), .RN(n1252), .Q(block[22]), 
        .QN(n381) );
  DFFRX1 \block_reg[38]  ( .D(n772), .CK(n1313), .RN(n1252), .Q(block[38]), 
        .QN(n380) );
  DFFRX1 \block_reg[54]  ( .D(n771), .CK(n1314), .RN(n1252), .Q(block[54]), 
        .QN(n379) );
  DFFRX1 \block_reg[70]  ( .D(n770), .CK(n1315), .RN(n1262), .Q(block[70]), 
        .QN(n378) );
  DFFRX1 \block_reg[86]  ( .D(n769), .CK(n1316), .RN(n1263), .Q(block[86]), 
        .QN(n377) );
  DFFRX1 \block_reg[102]  ( .D(n768), .CK(n1302), .RN(n1261), .Q(block[102]), 
        .QN(n376) );
  DFFRX1 \block_reg[118]  ( .D(n767), .CK(n1302), .RN(n1263), .Q(block[118]), 
        .QN(n375) );
  DFFRX1 \block_reg[111]  ( .D(n732), .CK(n1312), .RN(n1253), .Q(block[111]), 
        .QN(n341) );
  DFFRX1 \block_reg[79]  ( .D(n730), .CK(n1313), .RN(n1254), .Q(block[79]), 
        .QN(n339) );
  DFFRX1 \block_reg[47]  ( .D(n728), .CK(n1313), .RN(n1254), .Q(block[47]), 
        .QN(n337) );
  DFFRX1 \block_reg[15]  ( .D(n726), .CK(n1314), .RN(n1254), .Q(block[15]), 
        .QN(n335) );
  DFFRX1 \block_reg[7]  ( .D(n725), .CK(n1315), .RN(n1254), .Q(block[7]), .QN(
        n334) );
  DFFRX1 \block_reg[23]  ( .D(n724), .CK(n1316), .RN(n1254), .Q(block[23]), 
        .QN(n333) );
  DFFRX1 \block_reg[39]  ( .D(n723), .CK(n1310), .RN(n1254), .Q(block[39]), 
        .QN(n332) );
  DFFRX1 \block_reg[55]  ( .D(n722), .CK(n1308), .RN(n1254), .Q(block[55]), 
        .QN(n331) );
  DFFRX1 \block_reg[71]  ( .D(n721), .CK(n1312), .RN(n1254), .Q(block[71]), 
        .QN(n330) );
  DFFRX1 \block_reg[87]  ( .D(n720), .CK(n1308), .RN(n1255), .Q(block[87]), 
        .QN(n329) );
  DFFRX1 \block_reg[103]  ( .D(n719), .CK(n1315), .RN(n1255), .Q(block[103]), 
        .QN(n328) );
  DFFRX1 \block_reg[119]  ( .D(n718), .CK(n1304), .RN(n1255), .Q(block[119]), 
        .QN(n327) );
  DFFRX1 \key_reg[41]  ( .D(n1073), .CK(n1274), .RN(n1266), .Q(key[41]), .QN(
        n675) );
  DFFRX1 \key_reg[73]  ( .D(n1056), .CK(n1276), .RN(n1259), .Q(key[73]), .QN(
        n658) );
  DFFRX1 \key_reg[9]  ( .D(n1055), .CK(n1276), .RN(n1267), .Q(key[9]), .QN(
        n657) );
  DFFRX1 \key_reg[49]  ( .D(n1043), .CK(n1277), .RN(n1263), .Q(key[49]), .QN(
        n645) );
  DFFRX1 \key_reg[81]  ( .D(n1038), .CK(n1278), .RN(n1228), .Q(key[81]), .QN(
        n640) );
  DFFRX1 \key_reg[17]  ( .D(n1037), .CK(n1278), .RN(n1228), .Q(key[17]), .QN(
        n639) );
  DFFRX1 \key_reg[72]  ( .D(n1001), .CK(n1281), .RN(n1231), .Q(key[72]), .QN(
        n604) );
  DFFRX1 \key_reg[40]  ( .D(n999), .CK(n1281), .RN(n1232), .Q(key[40]), .QN(
        n602) );
  DFFRX1 \key_reg[8]  ( .D(n997), .CK(n1282), .RN(n1232), .Q(key[8]), .QN(n600) );
  DFFRX1 \key_reg[16]  ( .D(n995), .CK(n1282), .RN(n1232), .Q(key[16]), .QN(
        n598) );
  DFFRX1 \key_reg[48]  ( .D(n993), .CK(n1282), .RN(n1232), .Q(key[48]), .QN(
        n596) );
  DFFRX1 \key_reg[80]  ( .D(n991), .CK(n1282), .RN(n1232), .Q(key[80]), .QN(
        n594) );
  DFFRX1 \key_reg[76]  ( .D(n853), .CK(n1296), .RN(n1246), .Q(key[76]), .QN(
        n459) );
  DFFRX1 \key_reg[44]  ( .D(n851), .CK(n1296), .RN(n1246), .Q(key[44]), .QN(
        n457) );
  DFFRX1 \key_reg[20]  ( .D(n847), .CK(n1297), .RN(n1247), .Q(key[20]), .QN(
        n453) );
  DFFRX1 \key_reg[52]  ( .D(n845), .CK(n1297), .RN(n1247), .Q(key[52]), .QN(
        n451) );
  DFFRX1 \key_reg[46]  ( .D(n753), .CK(n1304), .RN(n1261), .Q(key[46]), .QN(
        n361) );
  DFFRX1 \key_reg[14]  ( .D(n751), .CK(clock), .RN(n1264), .Q(key[14]), .QN(
        n359) );
  DFFRX1 \key_reg[22]  ( .D(n749), .CK(n1312), .RN(n1259), .Q(key[22]), .QN(
        n357) );
  DFFRX1 \key_reg[86]  ( .D(n745), .CK(clock), .RN(n1260), .Q(key[86]), .QN(
        n353) );
  DFFRX1 \key_reg[233]  ( .D(n1076), .CK(n1274), .RN(n1265), .Q(key[233]), 
        .QN(n678) );
  DFFRX1 \key_reg[169]  ( .D(n1075), .CK(n1274), .RN(n1264), .Q(key[169]), 
        .QN(n677) );
  DFFRX1 \key_reg[249]  ( .D(n1070), .CK(n1274), .RN(n1263), .Q(key[249]), 
        .QN(n672) );
  DFFRX1 \key_reg[185]  ( .D(n1069), .CK(n1274), .RN(n1261), .Q(key[185]), 
        .QN(n671) );
  DFFRX1 \key_reg[217]  ( .D(n1064), .CK(n1275), .RN(n1266), .Q(key[217]), 
        .QN(n666) );
  DFFRX1 \key_reg[153]  ( .D(n1063), .CK(n1275), .RN(n1260), .Q(key[153]), 
        .QN(n665) );
  DFFRX1 \key_reg[201]  ( .D(n1058), .CK(n1276), .RN(n1266), .Q(key[201]), 
        .QN(n660) );
  DFFRX1 \key_reg[137]  ( .D(n1057), .CK(n1276), .RN(n1265), .Q(key[137]), 
        .QN(n659) );
  DFFRX1 \key_reg[225]  ( .D(n1052), .CK(n1276), .RN(n1262), .Q(key[225]), 
        .QN(n654) );
  DFFRX1 \key_reg[161]  ( .D(n1051), .CK(n1276), .RN(n1270), .Q(key[161]), 
        .QN(n653) );
  DFFRX1 \key_reg[241]  ( .D(n1046), .CK(n1277), .RN(n1260), .Q(key[241]), 
        .QN(n648) );
  DFFRX1 \key_reg[177]  ( .D(n1045), .CK(n1277), .RN(n1265), .Q(key[177]), 
        .QN(n647) );
  DFFRX1 \key_reg[209]  ( .D(n1040), .CK(n1277), .RN(n1228), .Q(key[209]), 
        .QN(n642) );
  DFFRX1 \key_reg[145]  ( .D(n1039), .CK(n1277), .RN(n1228), .Q(key[145]), 
        .QN(n641) );
  DFFRX1 \key_reg[193]  ( .D(n1034), .CK(n1278), .RN(n1228), .Q(key[193]), 
        .QN(n636) );
  DFFRX1 \key_reg[129]  ( .D(n1033), .CK(n1278), .RN(n1228), .Q(key[129]), 
        .QN(n635) );
  DFFRX1 \key_reg[248]  ( .D(n1012), .CK(n1280), .RN(n1230), .Q(key[248]), 
        .QN(n615) );
  DFFRX1 \key_reg[232]  ( .D(n1011), .CK(n1280), .RN(n1230), .Q(key[232]), 
        .QN(n614) );
  DFFRX1 \key_reg[216]  ( .D(n1010), .CK(n1280), .RN(n1231), .Q(key[216]), 
        .QN(n613) );
  DFFRX1 \key_reg[184]  ( .D(n1008), .CK(n1281), .RN(n1231), .Q(key[184]), 
        .QN(n611) );
  DFFRX1 \key_reg[152]  ( .D(n1006), .CK(n1281), .RN(n1231), .Q(key[152]), 
        .QN(n609) );
  DFFRX1 \key_reg[128]  ( .D(n988), .CK(n1283), .RN(n1233), .Q(key[128]), .QN(
        n591) );
  DFFRX1 \key_reg[144]  ( .D(n987), .CK(n1283), .RN(n1233), .Q(key[144]), .QN(
        n590) );
  DFFRX1 \key_reg[160]  ( .D(n986), .CK(n1283), .RN(n1233), .Q(key[160]), .QN(
        n589) );
  DFFRX1 \key_reg[176]  ( .D(n985), .CK(n1283), .RN(n1233), .Q(key[176]), .QN(
        n588) );
  DFFRX1 \key_reg[208]  ( .D(n983), .CK(n1283), .RN(n1233), .Q(key[208]), .QN(
        n586) );
  DFFRX1 \key_reg[224]  ( .D(n982), .CK(n1283), .RN(n1233), .Q(key[224]), .QN(
        n585) );
  DFFRX1 \key_reg[240]  ( .D(n981), .CK(n1283), .RN(n1233), .Q(key[240]), .QN(
        n584) );
  DFFRX1 \key_reg[250]  ( .D(n962), .CK(n1285), .RN(n1235), .Q(key[250]), .QN(
        n566) );
  DFFRX1 \key_reg[234]  ( .D(n961), .CK(n1285), .RN(n1235), .Q(key[234]), .QN(
        n565) );
  DFFRX1 \key_reg[218]  ( .D(n960), .CK(n1285), .RN(n1236), .Q(key[218]), .QN(
        n564) );
  DFFRX1 \key_reg[202]  ( .D(n959), .CK(n1285), .RN(n1236), .Q(key[202]), .QN(
        n563) );
  DFFRX1 \key_reg[186]  ( .D(n958), .CK(n1286), .RN(n1236), .Q(key[186]), .QN(
        n562) );
  DFFRX1 \key_reg[170]  ( .D(n957), .CK(n1286), .RN(n1236), .Q(key[170]), .QN(
        n561) );
  DFFRX1 \key_reg[154]  ( .D(n956), .CK(n1286), .RN(n1236), .Q(key[154]), .QN(
        n560) );
  DFFRX1 \key_reg[138]  ( .D(n955), .CK(n1286), .RN(n1236), .Q(key[138]), .QN(
        n559) );
  DFFRX1 \key_reg[130]  ( .D(n938), .CK(n1288), .RN(n1238), .Q(key[130]), .QN(
        n542) );
  DFFRX1 \key_reg[146]  ( .D(n937), .CK(n1288), .RN(n1238), .Q(key[146]), .QN(
        n541) );
  DFFRX1 \key_reg[162]  ( .D(n936), .CK(n1288), .RN(n1238), .Q(key[162]), .QN(
        n540) );
  DFFRX1 \key_reg[178]  ( .D(n935), .CK(n1288), .RN(n1238), .Q(key[178]), .QN(
        n539) );
  DFFRX1 \key_reg[194]  ( .D(n934), .CK(n1288), .RN(n1238), .Q(key[194]), .QN(
        n538) );
  DFFRX1 \key_reg[210]  ( .D(n933), .CK(n1288), .RN(n1238), .Q(key[210]), .QN(
        n537) );
  DFFRX1 \key_reg[226]  ( .D(n932), .CK(n1288), .RN(n1238), .Q(key[226]), .QN(
        n536) );
  DFFRX1 \key_reg[242]  ( .D(n931), .CK(n1288), .RN(n1238), .Q(key[242]), .QN(
        n535) );
  DFFRX1 \key_reg[251]  ( .D(n913), .CK(n1290), .RN(n1240), .Q(key[251]), .QN(
        n518) );
  DFFRX1 \key_reg[235]  ( .D(n912), .CK(n1290), .RN(n1240), .Q(key[235]), .QN(
        n517) );
  DFFRX1 \key_reg[219]  ( .D(n911), .CK(n1290), .RN(n1240), .Q(key[219]), .QN(
        n516) );
  DFFRX1 \key_reg[203]  ( .D(n910), .CK(n1290), .RN(n1241), .Q(key[203]), .QN(
        n515) );
  DFFRX1 \key_reg[187]  ( .D(n909), .CK(n1290), .RN(n1241), .Q(key[187]), .QN(
        n514) );
  DFFRX1 \key_reg[171]  ( .D(n908), .CK(n1291), .RN(n1241), .Q(key[171]), .QN(
        n513) );
  DFFRX1 \key_reg[155]  ( .D(n907), .CK(n1291), .RN(n1241), .Q(key[155]), .QN(
        n512) );
  DFFRX1 \key_reg[139]  ( .D(n906), .CK(n1291), .RN(n1241), .Q(key[139]), .QN(
        n511) );
  DFFRX1 \key_reg[131]  ( .D(n889), .CK(n1292), .RN(n1243), .Q(key[131]), .QN(
        n494) );
  DFFRX1 \key_reg[147]  ( .D(n888), .CK(n1293), .RN(n1243), .Q(key[147]), .QN(
        n493) );
  DFFRX1 \key_reg[163]  ( .D(n887), .CK(n1293), .RN(n1243), .Q(key[163]), .QN(
        n492) );
  DFFRX1 \key_reg[179]  ( .D(n886), .CK(n1293), .RN(n1243), .Q(key[179]), .QN(
        n491) );
  DFFRX1 \key_reg[195]  ( .D(n885), .CK(n1293), .RN(n1243), .Q(key[195]), .QN(
        n490) );
  DFFRX1 \key_reg[211]  ( .D(n884), .CK(n1293), .RN(n1243), .Q(key[211]), .QN(
        n489) );
  DFFRX1 \key_reg[227]  ( .D(n883), .CK(n1293), .RN(n1243), .Q(key[227]), .QN(
        n488) );
  DFFRX1 \key_reg[243]  ( .D(n882), .CK(n1293), .RN(n1243), .Q(key[243]), .QN(
        n487) );
  DFFRX1 \key_reg[252]  ( .D(n864), .CK(n1295), .RN(n1245), .Q(key[252]), .QN(
        n470) );
  DFFRX1 \key_reg[220]  ( .D(n862), .CK(n1295), .RN(n1245), .Q(key[220]), .QN(
        n468) );
  DFFRX1 \key_reg[204]  ( .D(n861), .CK(n1295), .RN(n1245), .Q(key[204]), .QN(
        n467) );
  DFFRX1 \key_reg[188]  ( .D(n860), .CK(n1295), .RN(n1246), .Q(key[188]), .QN(
        n466) );
  DFFRX1 \key_reg[172]  ( .D(n859), .CK(n1295), .RN(n1246), .Q(key[172]), .QN(
        n465) );
  DFFRX1 \key_reg[156]  ( .D(n858), .CK(n1296), .RN(n1246), .Q(key[156]), .QN(
        n464) );
  DFFRX1 \key_reg[140]  ( .D(n857), .CK(n1296), .RN(n1246), .Q(key[140]), .QN(
        n463) );
  DFFRX1 \key_reg[148]  ( .D(n839), .CK(n1297), .RN(n1269), .Q(key[148]), .QN(
        n445) );
  DFFRX1 \key_reg[164]  ( .D(n838), .CK(n1298), .RN(n1259), .Q(key[164]), .QN(
        n444) );
  DFFRX1 \key_reg[180]  ( .D(n837), .CK(n1298), .RN(n1260), .Q(key[180]), .QN(
        n443) );
  DFFRX1 \key_reg[212]  ( .D(n835), .CK(n1298), .RN(n1272), .Q(key[212]), .QN(
        n441) );
  DFFRX1 \key_reg[228]  ( .D(n834), .CK(n1298), .RN(n1267), .Q(key[228]), .QN(
        n440) );
  DFFRX1 \key_reg[244]  ( .D(n833), .CK(n1298), .RN(n1266), .Q(key[244]), .QN(
        n439) );
  DFFRX1 \key_reg[253]  ( .D(n815), .CK(n1300), .RN(n1248), .Q(key[253]), .QN(
        n422) );
  DFFRX1 \key_reg[237]  ( .D(n814), .CK(n1300), .RN(n1248), .Q(key[237]), .QN(
        n421) );
  DFFRX1 \key_reg[221]  ( .D(n813), .CK(n1300), .RN(n1248), .Q(key[221]), .QN(
        n420) );
  DFFRX1 \key_reg[205]  ( .D(n812), .CK(n1300), .RN(n1248), .Q(key[205]), .QN(
        n419) );
  DFFRX1 \key_reg[189]  ( .D(n811), .CK(n1300), .RN(n1248), .Q(key[189]), .QN(
        n418) );
  DFFRX1 \key_reg[173]  ( .D(n810), .CK(n1300), .RN(n1249), .Q(key[173]), .QN(
        n417) );
  DFFRX1 \key_reg[157]  ( .D(n809), .CK(n1300), .RN(n1249), .Q(key[157]), .QN(
        n416) );
  DFFRX1 \key_reg[141]  ( .D(n808), .CK(n1301), .RN(n1249), .Q(key[141]), .QN(
        n415) );
  DFFRX1 \key_reg[133]  ( .D(n791), .CK(n1306), .RN(n1250), .Q(key[133]), .QN(
        n398) );
  DFFRX1 \key_reg[149]  ( .D(n790), .CK(n1305), .RN(n1251), .Q(key[149]), .QN(
        n397) );
  DFFRX1 \key_reg[165]  ( .D(n789), .CK(n1303), .RN(n1251), .Q(key[165]), .QN(
        n396) );
  DFFRX1 \key_reg[181]  ( .D(n788), .CK(n1309), .RN(n1251), .Q(key[181]), .QN(
        n395) );
  DFFRX1 \key_reg[197]  ( .D(n787), .CK(n1308), .RN(n1251), .Q(key[197]), .QN(
        n394) );
  DFFRX1 \key_reg[213]  ( .D(n786), .CK(n1307), .RN(n1251), .Q(key[213]), .QN(
        n393) );
  DFFRX1 \key_reg[229]  ( .D(n785), .CK(n1304), .RN(n1251), .Q(key[229]), .QN(
        n392) );
  DFFRX1 \key_reg[245]  ( .D(n784), .CK(n1316), .RN(n1251), .Q(key[245]), .QN(
        n391) );
  DFFRX1 \key_reg[254]  ( .D(n766), .CK(n1302), .RN(n1260), .Q(key[254]), .QN(
        n374) );
  DFFRX1 \key_reg[238]  ( .D(n765), .CK(n1302), .RN(n1269), .Q(key[238]), .QN(
        n373) );
  DFFRX1 \key_reg[222]  ( .D(n764), .CK(n1302), .RN(n1271), .Q(key[222]), .QN(
        n372) );
  DFFRX1 \key_reg[190]  ( .D(n762), .CK(n1302), .RN(n1272), .Q(key[190]), .QN(
        n370) );
  DFFRX1 \key_reg[174]  ( .D(n761), .CK(n1302), .RN(n1268), .Q(key[174]), .QN(
        n369) );
  DFFRX1 \key_reg[158]  ( .D(n760), .CK(n1302), .RN(n1267), .Q(key[158]), .QN(
        n368) );
  DFFRX1 \key_reg[142]  ( .D(n759), .CK(n1302), .RN(n1266), .Q(key[142]), .QN(
        n367) );
  DFFRX1 \key_reg[134]  ( .D(n742), .CK(n1308), .RN(n1267), .Q(key[134]), .QN(
        n350) );
  DFFRX1 \key_reg[150]  ( .D(n741), .CK(n1306), .RN(n1266), .Q(key[150]), .QN(
        n349) );
  DFFRX1 \key_reg[166]  ( .D(n740), .CK(n1311), .RN(n1253), .Q(key[166]), .QN(
        n348) );
  DFFRX1 \key_reg[182]  ( .D(n739), .CK(n1310), .RN(n1253), .Q(key[182]), .QN(
        n347) );
  DFFRX1 \key_reg[198]  ( .D(n738), .CK(n1314), .RN(n1253), .Q(key[198]), .QN(
        n346) );
  DFFRX1 \key_reg[214]  ( .D(n737), .CK(n1315), .RN(n1253), .Q(key[214]), .QN(
        n345) );
  DFFRX1 \key_reg[230]  ( .D(n736), .CK(n1316), .RN(n1253), .Q(key[230]), .QN(
        n344) );
  DFFRX1 \key_reg[246]  ( .D(n735), .CK(n1306), .RN(n1253), .Q(key[246]), .QN(
        n343) );
  DFFRX1 \key_reg[255]  ( .D(n717), .CK(n1313), .RN(n1255), .Q(key[255]), .QN(
        n326) );
  DFFRX1 \key_reg[239]  ( .D(n716), .CK(n1308), .RN(n1255), .Q(key[239]), .QN(
        n325) );
  DFFRX1 \key_reg[223]  ( .D(n715), .CK(n1303), .RN(n1255), .Q(key[223]), .QN(
        n324) );
  DFFRX1 \key_reg[207]  ( .D(n714), .CK(n1303), .RN(n1255), .Q(key[207]), .QN(
        n323) );
  DFFRX1 \key_reg[191]  ( .D(n713), .CK(n1307), .RN(n1255), .Q(key[191]), .QN(
        n322) );
  DFFRX1 \key_reg[175]  ( .D(n712), .CK(n1311), .RN(n1255), .Q(key[175]), .QN(
        n321) );
  DFFRX1 \key_reg[159]  ( .D(n711), .CK(n1312), .RN(n1255), .Q(key[159]), .QN(
        n320) );
  DFFRX1 \key_reg[143]  ( .D(n710), .CK(n1310), .RN(n1256), .Q(key[143]), .QN(
        n319) );
  DFFRX1 \key_reg[135]  ( .D(n693), .CK(n1304), .RN(n1257), .Q(key[135]), .QN(
        n302) );
  DFFRX1 \key_reg[151]  ( .D(n692), .CK(n1314), .RN(n1257), .Q(key[151]), .QN(
        n301) );
  DFFRX1 \key_reg[167]  ( .D(n691), .CK(n1305), .RN(n1257), .Q(key[167]), .QN(
        n300) );
  DFFRX1 \key_reg[183]  ( .D(n690), .CK(n1303), .RN(n1258), .Q(key[183]), .QN(
        n299) );
  DFFRX1 \key_reg[199]  ( .D(n689), .CK(n1308), .RN(n1258), .Q(key[199]), .QN(
        n298) );
  DFFRX1 \key_reg[215]  ( .D(n688), .CK(n1306), .RN(n1258), .Q(key[215]), .QN(
        n297) );
  DFFRX1 \key_reg[231]  ( .D(n687), .CK(n1305), .RN(n1258), .Q(key[231]), .QN(
        n296) );
  DFFRX1 \key_reg[247]  ( .D(n686), .CK(n1310), .RN(n1258), .Q(key[247]), .QN(
        n295) );
  DFFRX1 \key_reg[105]  ( .D(n1074), .CK(n1274), .RN(n1263), .Q(key[105]), 
        .QN(n676) );
  DFFRX1 \key_reg[121]  ( .D(n1068), .CK(n1275), .RN(n1269), .Q(key[121]), 
        .QN(n670) );
  DFFRX1 \key_reg[57]  ( .D(n1067), .CK(n1275), .RN(n1270), .Q(key[57]), .QN(
        n669) );
  DFFRX1 \key_reg[89]  ( .D(n1062), .CK(n1275), .RN(n1272), .Q(key[89]), .QN(
        n664) );
  DFFRX1 \key_reg[25]  ( .D(n1061), .CK(n1275), .RN(n1271), .Q(key[25]), .QN(
        n663) );
  DFFRX1 \key_reg[97]  ( .D(n1050), .CK(n1276), .RN(n1269), .Q(key[97]), .QN(
        n652) );
  DFFRX1 \key_reg[33]  ( .D(n1049), .CK(n1276), .RN(n1270), .Q(key[33]), .QN(
        n651) );
  DFFRX1 \key_reg[113]  ( .D(n1044), .CK(n1277), .RN(n1269), .Q(key[113]), 
        .QN(n646) );
  DFFRX1 \key_reg[65]  ( .D(n1032), .CK(n1278), .RN(n1228), .Q(key[65]), .QN(
        n634) );
  DFFRX1 \key_reg[1]  ( .D(n1031), .CK(n1278), .RN(n1228), .Q(key[1]), .QN(
        n633) );
  DFFRX1 \key_reg[120]  ( .D(n1004), .CK(n1281), .RN(n1231), .Q(key[120]), 
        .QN(n607) );
  DFFRX1 \key_reg[104]  ( .D(n1003), .CK(n1281), .RN(n1231), .Q(key[104]), 
        .QN(n606) );
  DFFRX1 \key_reg[88]  ( .D(n1002), .CK(n1281), .RN(n1231), .Q(key[88]), .QN(
        n605) );
  DFFRX1 \key_reg[56]  ( .D(n1000), .CK(n1281), .RN(n1232), .Q(key[56]), .QN(
        n603) );
  DFFRX1 \key_reg[24]  ( .D(n998), .CK(n1282), .RN(n1232), .Q(key[24]), .QN(
        n601) );
  DFFRX1 \key_reg[0]  ( .D(n996), .CK(n1282), .RN(n1232), .Q(key[0]), .QN(n599) );
  DFFRX1 \key_reg[32]  ( .D(n994), .CK(n1282), .RN(n1232), .Q(key[32]), .QN(
        n597) );
  DFFRX1 \key_reg[64]  ( .D(n992), .CK(n1282), .RN(n1232), .Q(key[64]), .QN(
        n595) );
  DFFRX1 \key_reg[96]  ( .D(n990), .CK(n1282), .RN(n1233), .Q(key[96]), .QN(
        n593) );
  DFFRX1 \key_reg[112]  ( .D(n989), .CK(n1282), .RN(n1233), .Q(key[112]), .QN(
        n592) );
  DFFRX1 \key_reg[122]  ( .D(n954), .CK(n1286), .RN(n1236), .Q(key[122]), .QN(
        n558) );
  DFFRX1 \key_reg[106]  ( .D(n953), .CK(n1286), .RN(n1236), .Q(key[106]), .QN(
        n557) );
  DFFRX1 \key_reg[90]  ( .D(n952), .CK(n1286), .RN(n1236), .Q(key[90]), .QN(
        n556) );
  DFFRX1 \key_reg[74]  ( .D(n951), .CK(n1286), .RN(n1236), .Q(key[74]), .QN(
        n555) );
  DFFRX1 \key_reg[58]  ( .D(n950), .CK(n1286), .RN(n1237), .Q(key[58]), .QN(
        n554) );
  DFFRX1 \key_reg[42]  ( .D(n949), .CK(n1286), .RN(n1237), .Q(key[42]), .QN(
        n553) );
  DFFRX1 \key_reg[26]  ( .D(n948), .CK(n1287), .RN(n1237), .Q(key[26]), .QN(
        n552) );
  DFFRX1 \key_reg[10]  ( .D(n947), .CK(n1287), .RN(n1237), .Q(key[10]), .QN(
        n551) );
  DFFRX1 \key_reg[2]  ( .D(n946), .CK(n1287), .RN(n1237), .Q(key[2]), .QN(n550) );
  DFFRX1 \key_reg[18]  ( .D(n945), .CK(n1287), .RN(n1237), .Q(key[18]), .QN(
        n549) );
  DFFRX1 \key_reg[34]  ( .D(n944), .CK(n1287), .RN(n1237), .Q(key[34]), .QN(
        n548) );
  DFFRX1 \key_reg[50]  ( .D(n943), .CK(n1287), .RN(n1237), .Q(key[50]), .QN(
        n547) );
  DFFRX1 \key_reg[66]  ( .D(n942), .CK(n1287), .RN(n1237), .Q(key[66]), .QN(
        n546) );
  DFFRX1 \key_reg[82]  ( .D(n941), .CK(n1287), .RN(n1237), .Q(key[82]), .QN(
        n545) );
  DFFRX1 \key_reg[98]  ( .D(n940), .CK(n1287), .RN(n1238), .Q(key[98]), .QN(
        n544) );
  DFFRX1 \key_reg[114]  ( .D(n939), .CK(n1287), .RN(n1238), .Q(key[114]), .QN(
        n543) );
  DFFRX1 \key_reg[123]  ( .D(n905), .CK(n1291), .RN(n1241), .Q(key[123]), .QN(
        n510) );
  DFFRX1 \key_reg[107]  ( .D(n904), .CK(n1291), .RN(n1241), .Q(key[107]), .QN(
        n509) );
  DFFRX1 \key_reg[91]  ( .D(n903), .CK(n1291), .RN(n1241), .Q(key[91]), .QN(
        n508) );
  DFFRX1 \key_reg[75]  ( .D(n902), .CK(n1291), .RN(n1241), .Q(key[75]), .QN(
        n507) );
  DFFRX1 \key_reg[59]  ( .D(n901), .CK(n1291), .RN(n1241), .Q(key[59]), .QN(
        n506) );
  DFFRX1 \key_reg[43]  ( .D(n900), .CK(n1291), .RN(n1242), .Q(key[43]), .QN(
        n505) );
  DFFRX1 \key_reg[27]  ( .D(n899), .CK(n1291), .RN(n1242), .Q(key[27]), .QN(
        n504) );
  DFFRX1 \key_reg[11]  ( .D(n898), .CK(n1292), .RN(n1242), .Q(key[11]), .QN(
        n503) );
  DFFRX1 \key_reg[3]  ( .D(n897), .CK(n1292), .RN(n1242), .Q(key[3]), .QN(n502) );
  DFFRX1 \key_reg[19]  ( .D(n896), .CK(n1292), .RN(n1242), .Q(key[19]), .QN(
        n501) );
  DFFRX1 \key_reg[35]  ( .D(n895), .CK(n1292), .RN(n1242), .Q(key[35]), .QN(
        n500) );
  DFFRX1 \key_reg[51]  ( .D(n894), .CK(n1292), .RN(n1242), .Q(key[51]), .QN(
        n499) );
  DFFRX1 \key_reg[67]  ( .D(n893), .CK(n1292), .RN(n1242), .Q(key[67]), .QN(
        n498) );
  DFFRX1 \key_reg[83]  ( .D(n892), .CK(n1292), .RN(n1242), .Q(key[83]), .QN(
        n497) );
  DFFRX1 \key_reg[99]  ( .D(n891), .CK(n1292), .RN(n1242), .Q(key[99]), .QN(
        n496) );
  DFFRX1 \key_reg[115]  ( .D(n890), .CK(n1292), .RN(n1243), .Q(key[115]), .QN(
        n495) );
  DFFRX1 \key_reg[124]  ( .D(n856), .CK(n1296), .RN(n1246), .Q(key[124]), .QN(
        n462) );
  DFFRX1 \key_reg[108]  ( .D(n855), .CK(n1296), .RN(n1246), .Q(key[108]), .QN(
        n461) );
  DFFRX1 \key_reg[92]  ( .D(n854), .CK(n1296), .RN(n1246), .Q(key[92]), .QN(
        n460) );
  DFFRX1 \key_reg[60]  ( .D(n852), .CK(n1296), .RN(n1246), .Q(key[60]), .QN(
        n458) );
  DFFRX1 \key_reg[28]  ( .D(n850), .CK(n1296), .RN(n1247), .Q(key[28]), .QN(
        n456) );
  DFFRX1 \key_reg[4]  ( .D(n848), .CK(n1297), .RN(n1247), .Q(key[4]), .QN(n454) );
  DFFRX1 \key_reg[36]  ( .D(n846), .CK(n1297), .RN(n1247), .Q(key[36]), .QN(
        n452) );
  DFFRX1 \key_reg[68]  ( .D(n844), .CK(n1297), .RN(n1247), .Q(key[68]), .QN(
        n450) );
  DFFRX1 \key_reg[100]  ( .D(n842), .CK(n1297), .RN(n1247), .Q(key[100]), .QN(
        n448) );
  DFFRX1 \key_reg[116]  ( .D(n841), .CK(n1297), .RN(n1247), .Q(key[116]), .QN(
        n447) );
  DFFRX1 \key_reg[125]  ( .D(n807), .CK(n1301), .RN(n1249), .Q(key[125]), .QN(
        n414) );
  DFFRX1 \key_reg[109]  ( .D(n806), .CK(n1301), .RN(n1249), .Q(key[109]), .QN(
        n413) );
  DFFRX1 \key_reg[93]  ( .D(n805), .CK(n1301), .RN(n1249), .Q(key[93]), .QN(
        n412) );
  DFFRX1 \key_reg[77]  ( .D(n804), .CK(n1301), .RN(n1249), .Q(key[77]), .QN(
        n411) );
  DFFRX1 \key_reg[61]  ( .D(n803), .CK(n1301), .RN(n1249), .Q(key[61]), .QN(
        n410) );
  DFFRX1 \key_reg[45]  ( .D(n802), .CK(n1301), .RN(n1249), .Q(key[45]), .QN(
        n409) );
  DFFRX1 \key_reg[29]  ( .D(n801), .CK(n1301), .RN(n1249), .Q(key[29]), .QN(
        n408) );
  DFFRX1 \key_reg[13]  ( .D(n800), .CK(n1301), .RN(n1250), .Q(key[13]), .QN(
        n407) );
  DFFRX1 \key_reg[5]  ( .D(n799), .CK(n1301), .RN(n1250), .Q(key[5]), .QN(n406) );
  DFFRX1 \key_reg[21]  ( .D(n798), .CK(n1312), .RN(n1250), .Q(key[21]), .QN(
        n405) );
  DFFRX1 \key_reg[37]  ( .D(n797), .CK(n1313), .RN(n1250), .Q(key[37]), .QN(
        n404) );
  DFFRX1 \key_reg[53]  ( .D(n796), .CK(n1314), .RN(n1250), .Q(key[53]), .QN(
        n403) );
  DFFRX1 \key_reg[69]  ( .D(n795), .CK(n1315), .RN(n1250), .Q(key[69]), .QN(
        n402) );
  DFFRX1 \key_reg[85]  ( .D(n794), .CK(n1305), .RN(n1250), .Q(key[85]), .QN(
        n401) );
  DFFRX1 \key_reg[101]  ( .D(n793), .CK(n1316), .RN(n1250), .Q(key[101]), .QN(
        n400) );
  DFFRX1 \key_reg[117]  ( .D(n792), .CK(n1303), .RN(n1250), .Q(key[117]), .QN(
        n399) );
  DFFRX1 \key_reg[126]  ( .D(n758), .CK(n1313), .RN(n1272), .Q(key[126]), .QN(
        n366) );
  DFFRX1 \key_reg[110]  ( .D(n757), .CK(n1314), .RN(n1268), .Q(key[110]), .QN(
        n365) );
  DFFRX1 \key_reg[94]  ( .D(n756), .CK(n1303), .RN(n1269), .Q(key[94]), .QN(
        n364) );
  DFFRX1 \key_reg[62]  ( .D(n754), .CK(n1316), .RN(n1270), .Q(key[62]), .QN(
        n362) );
  DFFRX1 \key_reg[30]  ( .D(n752), .CK(n1308), .RN(n1271), .Q(key[30]), .QN(
        n360) );
  DFFRX1 \key_reg[6]  ( .D(n750), .CK(n1303), .RN(n1265), .Q(key[6]), .QN(n358) );
  DFFRX1 \key_reg[38]  ( .D(n748), .CK(n1309), .RN(n1264), .Q(key[38]), .QN(
        n356) );
  DFFRX1 \key_reg[70]  ( .D(n746), .CK(n1315), .RN(n1263), .Q(key[70]), .QN(
        n354) );
  DFFRX1 \key_reg[102]  ( .D(n744), .CK(n1305), .RN(n1262), .Q(key[102]), .QN(
        n352) );
  DFFRX1 \key_reg[118]  ( .D(n743), .CK(n1303), .RN(n1265), .Q(key[118]), .QN(
        n351) );
  DFFRX1 \key_reg[127]  ( .D(n709), .CK(n1311), .RN(n1256), .Q(key[127]), .QN(
        n318) );
  DFFRX1 \key_reg[111]  ( .D(n708), .CK(n1314), .RN(n1256), .Q(key[111]), .QN(
        n317) );
  DFFRX1 \key_reg[95]  ( .D(n707), .CK(n1309), .RN(n1256), .Q(key[95]), .QN(
        n316) );
  DFFRX1 \key_reg[79]  ( .D(n706), .CK(n1316), .RN(n1256), .Q(key[79]), .QN(
        n315) );
  DFFRX1 \key_reg[63]  ( .D(n705), .CK(n1307), .RN(n1256), .Q(key[63]), .QN(
        n314) );
  DFFRX1 \key_reg[47]  ( .D(n704), .CK(n1315), .RN(n1256), .Q(key[47]), .QN(
        n313) );
  DFFRX1 \key_reg[31]  ( .D(n703), .CK(n1309), .RN(n1256), .Q(key[31]), .QN(
        n312) );
  DFFRX1 \key_reg[15]  ( .D(n702), .CK(n1311), .RN(n1256), .Q(key[15]), .QN(
        n311) );
  DFFRX1 \key_reg[7]  ( .D(n701), .CK(n1310), .RN(n1256), .Q(key[7]), .QN(n310) );
  DFFRX1 \key_reg[23]  ( .D(n700), .CK(n1312), .RN(n1257), .Q(key[23]), .QN(
        n309) );
  DFFRX1 \key_reg[39]  ( .D(n699), .CK(n1313), .RN(n1257), .Q(key[39]), .QN(
        n308) );
  DFFRX1 \key_reg[55]  ( .D(n698), .CK(n1314), .RN(n1257), .Q(key[55]), .QN(
        n307) );
  DFFRX1 \key_reg[71]  ( .D(n697), .CK(n1312), .RN(n1257), .Q(key[71]), .QN(
        n306) );
  DFFRX1 \key_reg[87]  ( .D(n696), .CK(n1313), .RN(n1257), .Q(key[87]), .QN(
        n305) );
  DFFRX1 \key_reg[103]  ( .D(n695), .CK(n1307), .RN(n1257), .Q(key[103]), .QN(
        n304) );
  DFFRX1 \key_reg[119]  ( .D(n694), .CK(n1306), .RN(n1257), .Q(key[119]), .QN(
        n303) );
  DFFRX1 \key_reg[200]  ( .D(n1009), .CK(n1280), .RN(n1231), .Q(key[200]), 
        .QN(n612) );
  DFFRX1 \key_reg[168]  ( .D(n1007), .CK(n1281), .RN(n1231), .Q(key[168]), 
        .QN(n610) );
  DFFRX1 \key_reg[136]  ( .D(n1005), .CK(n1281), .RN(n1231), .Q(key[136]), 
        .QN(n608) );
  DFFRX1 \key_reg[192]  ( .D(n984), .CK(n1283), .RN(n1233), .Q(key[192]), .QN(
        n587) );
  DFFRX1 \key_reg[236]  ( .D(n863), .CK(n1295), .RN(n1245), .Q(key[236]), .QN(
        n469) );
  DFFRX1 \key_reg[132]  ( .D(n840), .CK(n1297), .RN(n1265), .Q(key[132]), .QN(
        n446) );
  DFFRX1 \key_reg[196]  ( .D(n836), .CK(n1298), .RN(n1262), .Q(key[196]), .QN(
        n442) );
  DFFRX1 \key_reg[206]  ( .D(n763), .CK(n1302), .RN(n1264), .Q(key[206]), .QN(
        n371) );
  DFFRX1 \key_reg[12]  ( .D(n849), .CK(n1296), .RN(n1247), .Q(key[12]), .QN(
        n455) );
  DFFRX1 \key_reg[84]  ( .D(n843), .CK(n1297), .RN(n1247), .Q(key[84]), .QN(
        n449) );
  DFFRX1 \next_status_reg[1]  ( .D(n1082), .CK(n1273), .RN(n1272), .Q(
        next_status[1]), .QN(n1096) );
  DFFRX1 encdec_reg ( .D(n980), .CK(n1283), .RN(n1234), .Q(encdec), .QN(n583)
         );
  DFFRX1 \block_reg[57]  ( .D(n1066), .CK(n1275), .RN(n1262), .Q(block[57]), 
        .QN(n668) );
  DFFRX1 \block_reg[121]  ( .D(n1065), .CK(n1275), .RN(n1259), .Q(block[121]), 
        .QN(n667) );
  DFFRX1 \block_reg[25]  ( .D(n1060), .CK(n1275), .RN(n1264), .Q(block[25]), 
        .QN(n662) );
  DFFRX1 \block_reg[89]  ( .D(n1059), .CK(n1275), .RN(n1261), .Q(block[89]), 
        .QN(n661) );
  DFFRX1 \block_reg[120]  ( .D(n1027), .CK(n1279), .RN(n1229), .Q(block[120]), 
        .QN(n630) );
  DFFRX1 \block_reg[88]  ( .D(n1025), .CK(n1279), .RN(n1229), .Q(block[88]), 
        .QN(n628) );
  DFFRX1 \block_reg[56]  ( .D(n1023), .CK(n1279), .RN(n1229), .Q(block[56]), 
        .QN(n626) );
  DFFRX1 \block_reg[24]  ( .D(n1021), .CK(n1279), .RN(n1229), .Q(block[24]), 
        .QN(n624) );
  DFFRX1 \block_reg[122]  ( .D(n978), .CK(n1284), .RN(n1234), .Q(block[122]), 
        .QN(n582) );
  DFFRX1 \block_reg[90]  ( .D(n976), .CK(n1284), .RN(n1234), .Q(block[90]), 
        .QN(n580) );
  DFFRX1 \block_reg[58]  ( .D(n974), .CK(n1284), .RN(n1234), .Q(block[58]), 
        .QN(n578) );
  DFFRX1 \block_reg[26]  ( .D(n972), .CK(n1284), .RN(n1234), .Q(block[26]), 
        .QN(n576) );
  DFFRX1 \block_reg[123]  ( .D(n929), .CK(n1288), .RN(n1239), .Q(block[123]), 
        .QN(n534) );
  DFFRX1 \block_reg[91]  ( .D(n927), .CK(n1289), .RN(n1239), .Q(block[91]), 
        .QN(n532) );
  DFFRX1 \block_reg[59]  ( .D(n925), .CK(n1289), .RN(n1239), .Q(block[59]), 
        .QN(n530) );
  DFFRX1 \block_reg[27]  ( .D(n923), .CK(n1289), .RN(n1239), .Q(block[27]), 
        .QN(n528) );
  DFFRX1 \block_reg[124]  ( .D(n880), .CK(n1293), .RN(n1244), .Q(block[124]), 
        .QN(n486) );
  DFFRX1 \block_reg[92]  ( .D(n878), .CK(n1294), .RN(n1244), .Q(block[92]), 
        .QN(n484) );
  DFFRX1 \block_reg[60]  ( .D(n876), .CK(n1294), .RN(n1244), .Q(block[60]), 
        .QN(n482) );
  DFFRX1 \block_reg[28]  ( .D(n874), .CK(n1294), .RN(n1244), .Q(block[28]), 
        .QN(n480) );
  DFFRX1 \block_reg[125]  ( .D(n831), .CK(n1298), .RN(n1270), .Q(block[125]), 
        .QN(n438) );
  DFFRX1 \block_reg[93]  ( .D(n829), .CK(n1298), .RN(n1260), .Q(block[93]), 
        .QN(n436) );
  DFFRX1 \block_reg[61]  ( .D(n827), .CK(n1299), .RN(n1272), .Q(block[61]), 
        .QN(n434) );
  DFFRX1 \block_reg[29]  ( .D(n825), .CK(n1299), .RN(n1261), .Q(block[29]), 
        .QN(n432) );
  DFFRX1 \block_reg[126]  ( .D(n782), .CK(n1303), .RN(n1251), .Q(block[126]), 
        .QN(n390) );
  DFFRX1 \block_reg[94]  ( .D(n780), .CK(n1306), .RN(n1252), .Q(block[94]), 
        .QN(n388) );
  DFFRX1 \block_reg[62]  ( .D(n778), .CK(n1310), .RN(n1252), .Q(block[62]), 
        .QN(n386) );
  DFFRX1 \block_reg[30]  ( .D(n776), .CK(n1309), .RN(n1252), .Q(block[30]), 
        .QN(n384) );
  DFFRX1 \block_reg[127]  ( .D(n733), .CK(n1309), .RN(n1253), .Q(block[127]), 
        .QN(n342) );
  DFFRX1 \block_reg[95]  ( .D(n731), .CK(n1311), .RN(n1253), .Q(block[95]), 
        .QN(n340) );
  DFFRX1 \block_reg[63]  ( .D(n729), .CK(n1304), .RN(n1254), .Q(block[63]), 
        .QN(n338) );
  DFFRX1 \block_reg[31]  ( .D(n727), .CK(n1316), .RN(n1254), .Q(block[31]), 
        .QN(n336) );
  DFFRX1 \next_status_reg[2]  ( .D(n1083), .CK(n1273), .RN(n1268), .Q(
        next_status[2]), .QN(n1154) );
  DFFRX1 \next_status_reg[0]  ( .D(n1081), .CK(n1273), .RN(n1269), .Q(
        next_status[0]), .QN(n1101) );
  DFFRX1 next_reg ( .D(N58), .CK(sysclock), .RN(n1258), .Q(next) );
  DFFRX1 \current_status_reg[1]  ( .D(next_status[1]), .CK(sysclock), .RN(
        n1258), .Q(phase[1]) );
  DFFRX1 init_reg ( .D(N57), .CK(sysclock), .RN(n1258), .Q(init) );
  DFFRX1 \cnt_32_reg[4]  ( .D(n1084), .CK(n1273), .RN(n1270), .Q(cnt_32[4]), 
        .QN(n684) );
  DFFRX1 \cnt_32_reg[2]  ( .D(n1078), .CK(n1274), .RN(n1262), .Q(cnt_32[2]), 
        .QN(n680) );
  DFFRX1 \cnt_32_reg[1]  ( .D(n1079), .CK(n1273), .RN(n1265), .Q(cnt_32[1]), 
        .QN(n681) );
  DFFRX1 \cnt_32_reg[0]  ( .D(n1085), .CK(n1273), .RN(n1271), .Q(cnt_32[0]), 
        .QN(n682) );
  DFFRX1 \result_reg_reg[1]  ( .D(n1087), .CK(n1273), .RN(n1267), .Q(
        result_reg[1]), .QN(n1099) );
  DFFRX1 \result_reg_reg[0]  ( .D(n1028), .CK(n1279), .RN(n1229), .Q(
        result_reg[0]), .QN(n1098) );
  DFFRX1 \result_reg_reg[2]  ( .D(n979), .CK(n1283), .RN(n1234), .Q(
        result_reg[2]), .QN(n1100) );
  DFFRX1 \result_reg_reg[3]  ( .D(n930), .CK(n1288), .RN(n1239), .Q(
        result_reg[3]), .QN(n1094) );
  DFFRX1 \result_reg_reg[4]  ( .D(n881), .CK(n1293), .RN(n1243), .Q(
        result_reg[4]), .QN(n1095) );
  DFFRX1 \result_reg_reg[5]  ( .D(n832), .CK(n1298), .RN(n1271), .Q(
        result_reg[5]), .QN(n1093) );
  DFFRX1 \result_reg_reg[6]  ( .D(n783), .CK(n1311), .RN(n1251), .Q(
        result_reg[6]), .QN(n1092) );
  DFFRX1 \result_reg_reg[7]  ( .D(n734), .CK(n1309), .RN(n1253), .Q(
        result_reg[7]), .QN(n1091) );
  DFFRX1 \current_status_reg[0]  ( .D(next_status[0]), .CK(sysclock), .RN(
        n1258), .Q(phase[0]) );
  DFFRX1 \current_status_reg[2]  ( .D(next_status[2]), .CK(sysclock), .RN(
        n1258), .Q(phase[2]), .QN(n1097) );
  DFFRX1 keylen_reg ( .D(n1086), .CK(n1273), .RN(n1263), .Q(keylen), .QN(n679)
         );
  DFFRX1 \cnt_32_reg[3]  ( .D(n1077), .CK(n1274), .RN(n1261), .Q(cnt_32[3]), 
        .QN(n683) );
  BUFX2 U706 ( .A(keylen), .Y(n1102) );
  OAI2BB1XL U707 ( .A0N(cnt_32[4]), .A1N(n1319), .B0(keylen), .Y(n1318) );
  INVX1 U708 ( .A(n137), .Y(n1322) );
  OAI22XL U709 ( .A0(n1191), .A1(n1099), .B0(n1326), .B1(n1090), .Y(
        display_data[1]) );
  INVX3 U710 ( .A(n1090), .Y(n1191) );
  NOR2X1 U711 ( .A(n131), .B(cnt_32[2]), .Y(n222) );
  OAI21XL U712 ( .A0(n232), .A1(n113), .B0(n132), .Y(n112) );
  NAND2X1 U713 ( .A(cnt_32[4]), .B(cnt_32[3]), .Y(n170) );
  OAI2BB2XL U714 ( .B0(n1189), .B1(n1100), .A0N(data[2]), .A1N(n1191), .Y(
        display_data[2]) );
  OAI2BB2XL U715 ( .B0(n1190), .B1(n1094), .A0N(data[3]), .A1N(n1089), .Y(
        display_data[3]) );
  OAI2BB2XL U716 ( .B0(n1191), .B1(n1092), .A0N(data[6]), .A1N(n1089), .Y(
        display_data[6]) );
  OAI2BB2XL U717 ( .B0(n1191), .B1(n1093), .A0N(data[5]), .A1N(n1089), .Y(
        display_data[5]) );
  OAI2BB2XL U718 ( .B0(n1191), .B1(n1091), .A0N(data[7]), .A1N(n1089), .Y(
        display_data[7]) );
  NAND3X1 U719 ( .A(phase[1]), .B(n1097), .C(phase[0]), .Y(n239) );
  NOR2X1 U720 ( .A(n131), .B(n680), .Y(n213) );
  NAND2X1 U721 ( .A(n683), .B(cnt_32[4]), .Y(n154) );
  NAND2X1 U722 ( .A(n684), .B(cnt_32[3]), .Y(n204) );
  NAND2X1 U723 ( .A(n684), .B(n683), .Y(n185) );
  NAND2X1 U724 ( .A(n681), .B(cnt_32[0]), .Y(n226) );
  NAND2X1 U725 ( .A(n681), .B(n682), .Y(n223) );
  BUFX2 U726 ( .A(n1322), .Y(n1184) );
  BUFX2 U727 ( .A(n1322), .Y(n1185) );
  BUFX2 U728 ( .A(n1322), .Y(n1187) );
  BUFX2 U729 ( .A(n1322), .Y(n1186) );
  BUFX2 U730 ( .A(n1322), .Y(n1188) );
  BUFX2 U731 ( .A(n1259), .Y(n1257) );
  BUFX2 U732 ( .A(n1259), .Y(n1256) );
  BUFX2 U733 ( .A(n1260), .Y(n1255) );
  BUFX2 U734 ( .A(n1260), .Y(n1254) );
  BUFX2 U735 ( .A(n1260), .Y(n1253) );
  BUFX2 U736 ( .A(n1271), .Y(n1252) );
  BUFX2 U737 ( .A(n1272), .Y(n1251) );
  BUFX2 U738 ( .A(n1270), .Y(n1250) );
  BUFX2 U739 ( .A(n1261), .Y(n1249) );
  BUFX2 U740 ( .A(n1261), .Y(n1248) );
  BUFX2 U741 ( .A(n1266), .Y(n1247) );
  BUFX2 U742 ( .A(n1267), .Y(n1246) );
  BUFX2 U743 ( .A(n1262), .Y(n1245) );
  BUFX2 U744 ( .A(n1262), .Y(n1244) );
  BUFX2 U745 ( .A(n1262), .Y(n1243) );
  BUFX2 U746 ( .A(n1263), .Y(n1242) );
  BUFX2 U747 ( .A(n1263), .Y(n1241) );
  BUFX2 U748 ( .A(n1263), .Y(n1240) );
  BUFX2 U749 ( .A(n1264), .Y(n1239) );
  BUFX2 U750 ( .A(n1264), .Y(n1238) );
  BUFX2 U751 ( .A(n1264), .Y(n1237) );
  BUFX2 U752 ( .A(n1265), .Y(n1236) );
  BUFX2 U753 ( .A(n1265), .Y(n1235) );
  BUFX2 U754 ( .A(n1265), .Y(n1234) );
  BUFX2 U755 ( .A(n1266), .Y(n1233) );
  BUFX2 U756 ( .A(n1266), .Y(n1232) );
  BUFX2 U757 ( .A(n1266), .Y(n1231) );
  BUFX2 U758 ( .A(n1267), .Y(n1230) );
  BUFX2 U759 ( .A(n1267), .Y(n1229) );
  BUFX2 U760 ( .A(n1267), .Y(n1228) );
  BUFX2 U761 ( .A(n1259), .Y(n1258) );
  BUFX2 U762 ( .A(n1321), .Y(n1181) );
  BUFX2 U763 ( .A(n1303), .Y(n1302) );
  BUFX2 U764 ( .A(clock), .Y(n1301) );
  BUFX2 U765 ( .A(n1304), .Y(n1300) );
  BUFX2 U766 ( .A(n1307), .Y(n1299) );
  BUFX2 U767 ( .A(n1304), .Y(n1298) );
  BUFX2 U768 ( .A(n1304), .Y(n1297) );
  BUFX2 U769 ( .A(n1304), .Y(n1296) );
  BUFX2 U770 ( .A(n1305), .Y(n1295) );
  BUFX2 U771 ( .A(n1305), .Y(n1294) );
  BUFX2 U772 ( .A(n1305), .Y(n1293) );
  BUFX2 U773 ( .A(n1306), .Y(n1292) );
  BUFX2 U774 ( .A(n1306), .Y(n1291) );
  BUFX2 U775 ( .A(n1306), .Y(n1290) );
  BUFX2 U776 ( .A(n1307), .Y(n1289) );
  BUFX2 U777 ( .A(n1307), .Y(n1288) );
  BUFX2 U778 ( .A(n1307), .Y(n1287) );
  BUFX2 U779 ( .A(n1308), .Y(n1286) );
  BUFX2 U780 ( .A(n1308), .Y(n1285) );
  BUFX2 U781 ( .A(n1308), .Y(n1284) );
  BUFX2 U782 ( .A(n1309), .Y(n1283) );
  BUFX2 U783 ( .A(n1309), .Y(n1282) );
  BUFX2 U784 ( .A(n1309), .Y(n1281) );
  BUFX2 U785 ( .A(n1310), .Y(n1280) );
  BUFX2 U786 ( .A(n1310), .Y(n1279) );
  BUFX2 U787 ( .A(n1310), .Y(n1278) );
  BUFX2 U788 ( .A(n1311), .Y(n1277) );
  BUFX2 U789 ( .A(n1311), .Y(n1276) );
  BUFX2 U790 ( .A(n1311), .Y(n1275) );
  BUFX2 U791 ( .A(n1312), .Y(n1274) );
  BUFX2 U792 ( .A(n1312), .Y(n1273) );
  NAND2X1 U793 ( .A(n112), .B(n113), .Y(n9) );
  OAI22XL U794 ( .A0(n1181), .A1(n113), .B0(n1191), .B1(n112), .Y(n1080) );
  NAND2X1 U795 ( .A(n238), .B(n1184), .Y(n235) );
  OAI21XL U796 ( .A0(n1183), .A1(n125), .B0(n1325), .Y(n238) );
  NAND2X1 U797 ( .A(n222), .B(n29), .Y(n180) );
  NAND2X1 U798 ( .A(n222), .B(n1327), .Y(n174) );
  NAND2X1 U799 ( .A(n222), .B(n1329), .Y(n171) );
  NAND2X1 U800 ( .A(n222), .B(n26), .Y(n177) );
  NAND2X1 U801 ( .A(n1182), .B(n1325), .Y(n131) );
  OA21XL U802 ( .A0(n170), .A1(n167), .B0(n1185), .Y(n1103) );
  INVX1 U803 ( .A(n1103), .Y(n160) );
  OA21XL U804 ( .A0(n170), .A1(n159), .B0(n1187), .Y(n1104) );
  INVX1 U805 ( .A(n1104), .Y(n188) );
  OA21XL U806 ( .A0(n170), .A1(n174), .B0(n1188), .Y(n1105) );
  INVX1 U807 ( .A(n1105), .Y(n172) );
  OA21XL U808 ( .A0(n170), .A1(n180), .B0(n1188), .Y(n1106) );
  INVX1 U809 ( .A(n1106), .Y(n178) );
  OA21XL U810 ( .A0(n164), .A1(n170), .B0(n1186), .Y(n1107) );
  INVX1 U811 ( .A(n1107), .Y(n140) );
  OA21XL U812 ( .A0(n170), .A1(n155), .B0(n1188), .Y(n1108) );
  INVX1 U813 ( .A(n1108), .Y(n181) );
  OA21XL U814 ( .A0(n1330), .A1(n269), .B0(n1184), .Y(n1109) );
  INVX1 U815 ( .A(n1109), .Y(n274) );
  OA21XL U816 ( .A0(n1328), .A1(n279), .B0(n1184), .Y(n1110) );
  INVX1 U817 ( .A(n1110), .Y(n241) );
  OA21XL U818 ( .A0(n170), .A1(n171), .B0(n1188), .Y(n1111) );
  INVX1 U819 ( .A(n1111), .Y(n168) );
  OA21XL U820 ( .A0(n1328), .A1(n269), .B0(n1185), .Y(n1112) );
  INVX1 U821 ( .A(n1112), .Y(n272) );
  OA21XL U822 ( .A0(n170), .A1(n177), .B0(n1188), .Y(n1113) );
  INVX1 U823 ( .A(n1113), .Y(n175) );
  OA21XL U824 ( .A0(n1330), .A1(n279), .B0(n1186), .Y(n1114) );
  INVX1 U825 ( .A(n1114), .Y(n258) );
  BUFX2 U826 ( .A(n19), .Y(n1222) );
  BUFX2 U827 ( .A(n18), .Y(n1225) );
  INVX1 U828 ( .A(n112), .Y(n1321) );
  INVX1 U829 ( .A(n129), .Y(n1182) );
  INVX1 U830 ( .A(n129), .Y(n1183) );
  BUFX2 U831 ( .A(n19), .Y(n1223) );
  BUFX2 U832 ( .A(n18), .Y(n1226) );
  BUFX2 U833 ( .A(n1272), .Y(n1260) );
  BUFX2 U834 ( .A(n1305), .Y(n1303) );
  BUFX2 U835 ( .A(n1271), .Y(n1261) );
  BUFX2 U836 ( .A(n1315), .Y(n1304) );
  BUFX2 U837 ( .A(n1316), .Y(n1305) );
  BUFX2 U838 ( .A(n1270), .Y(n1262) );
  BUFX2 U839 ( .A(n1316), .Y(n1306) );
  BUFX2 U840 ( .A(n1270), .Y(n1263) );
  BUFX2 U841 ( .A(n1315), .Y(n1307) );
  BUFX2 U842 ( .A(n1269), .Y(n1264) );
  BUFX2 U843 ( .A(n1315), .Y(n1308) );
  BUFX2 U844 ( .A(n1269), .Y(n1265) );
  BUFX2 U845 ( .A(n1314), .Y(n1309) );
  BUFX2 U846 ( .A(n1268), .Y(n1266) );
  BUFX2 U847 ( .A(n1314), .Y(n1310) );
  BUFX2 U848 ( .A(n1268), .Y(n1267) );
  BUFX2 U849 ( .A(n1313), .Y(n1311) );
  BUFX2 U850 ( .A(n1272), .Y(n1259) );
  INVX1 U851 ( .A(n26), .Y(n1328) );
  INVX1 U852 ( .A(n29), .Y(n1330) );
  BUFX2 U853 ( .A(n1313), .Y(n1312) );
  BUFX2 U854 ( .A(n18), .Y(n1227) );
  BUFX2 U855 ( .A(n19), .Y(n1224) );
  OAI22XL U856 ( .A0(n1191), .A1(n1098), .B0(n1332), .B1(n1090), .Y(
        display_data[0]) );
  INVX4 U857 ( .A(n1090), .Y(n1189) );
  INVX4 U858 ( .A(n1090), .Y(n1190) );
  OAI211X1 U859 ( .A0(N94), .A1(n131), .B0(n132), .C0(n133), .Y(n121) );
  AOI31X1 U860 ( .A0(n125), .A1(n1331), .A2(n1325), .B0(n1324), .Y(n133) );
  INVX1 U861 ( .A(N108), .Y(n1331) );
  NOR3X1 U862 ( .A(n1097), .B(n233), .C(n232), .Y(n137) );
  NAND2X1 U863 ( .A(n233), .B(n1097), .Y(n113) );
  NAND2X1 U864 ( .A(n116), .B(cnt_32[3]), .Y(n18) );
  NAND2X1 U865 ( .A(n117), .B(cnt_32[3]), .Y(n19) );
  NOR3X1 U866 ( .A(cnt_32[4]), .B(n232), .C(n239), .Y(n291) );
  NOR2X1 U867 ( .A(cnt_32[2]), .B(n1181), .Y(n117) );
  INVX1 U868 ( .A(n239), .Y(n1323) );
  NAND2X1 U869 ( .A(n213), .B(n26), .Y(n164) );
  NAND2X1 U870 ( .A(n276), .B(cnt_32[3]), .Y(n269) );
  NAND2X1 U871 ( .A(n266), .B(cnt_32[3]), .Y(n279) );
  NAND2X1 U872 ( .A(n213), .B(n29), .Y(n167) );
  NAND2X1 U873 ( .A(n213), .B(n1327), .Y(n159) );
  NAND2X1 U874 ( .A(n213), .B(n1329), .Y(n155) );
  NAND2X1 U875 ( .A(n239), .B(n113), .Y(n125) );
  OA21XL U876 ( .A0(n154), .A1(n167), .B0(n1188), .Y(n1115) );
  INVX1 U877 ( .A(n1115), .Y(n165) );
  OA21XL U878 ( .A0(n154), .A1(n159), .B0(n1188), .Y(n1116) );
  INVX1 U879 ( .A(n1116), .Y(n157) );
  OA21XL U880 ( .A0(n154), .A1(n174), .B0(n1186), .Y(n1117) );
  INVX1 U881 ( .A(n1117), .Y(n224) );
  OA21XL U882 ( .A0(n154), .A1(n155), .B0(n1184), .Y(n1118) );
  INVX1 U883 ( .A(n1118), .Y(n148) );
  OA21XL U884 ( .A0(n154), .A1(n171), .B0(n1186), .Y(n1119) );
  INVX1 U885 ( .A(n1119), .Y(n220) );
  OA21XL U886 ( .A0(n154), .A1(n177), .B0(n1185), .Y(n1120) );
  INVX1 U887 ( .A(n1120), .Y(n227) );
  OA21XL U888 ( .A0(n180), .A1(n154), .B0(n1185), .Y(n1121) );
  INVX1 U889 ( .A(n1121), .Y(n143) );
  OA21XL U890 ( .A0(n164), .A1(n154), .B0(n1188), .Y(n1122) );
  INVX1 U891 ( .A(n1122), .Y(n162) );
  OA21XL U892 ( .A0(n167), .A1(n185), .B0(n1187), .Y(n1123) );
  INVX1 U893 ( .A(n1123), .Y(n200) );
  OA21XL U894 ( .A0(n159), .A1(n185), .B0(n1187), .Y(n1124) );
  INVX1 U895 ( .A(n1124), .Y(n196) );
  OA21XL U896 ( .A0(n174), .A1(n185), .B0(n1187), .Y(n1125) );
  INVX1 U897 ( .A(n1125), .Y(n186) );
  OA21XL U898 ( .A0(n180), .A1(n185), .B0(n1187), .Y(n1126) );
  INVX1 U899 ( .A(n1126), .Y(n192) );
  OA21XL U900 ( .A0(n164), .A1(n185), .B0(n1187), .Y(n1127) );
  INVX1 U901 ( .A(n1127), .Y(n198) );
  OA21XL U902 ( .A0(n155), .A1(n185), .B0(n1187), .Y(n1128) );
  INVX1 U903 ( .A(n1128), .Y(n194) );
  OA21XL U904 ( .A0(n171), .A1(n185), .B0(n1188), .Y(n1129) );
  INVX1 U905 ( .A(n1129), .Y(n183) );
  OA21XL U906 ( .A0(n177), .A1(n185), .B0(n1187), .Y(n1130) );
  INVX1 U907 ( .A(n1130), .Y(n190) );
  OA21XL U908 ( .A0(n1330), .A1(n255), .B0(n1185), .Y(n1131) );
  INVX1 U909 ( .A(n1131), .Y(n263) );
  OA21XL U910 ( .A0(n167), .A1(n204), .B0(n1186), .Y(n1132) );
  INVX1 U911 ( .A(n1132), .Y(n218) );
  OA21XL U912 ( .A0(n226), .A1(n255), .B0(n1185), .Y(n1133) );
  INVX1 U913 ( .A(n1133), .Y(n256) );
  OA21XL U914 ( .A0(n226), .A1(n279), .B0(n1184), .Y(n1134) );
  INVX1 U915 ( .A(n1134), .Y(n280) );
  OA21XL U916 ( .A0(n159), .A1(n204), .B0(n1186), .Y(n1135) );
  INVX1 U917 ( .A(n1135), .Y(n214) );
  OA21XL U918 ( .A0(n226), .A1(n284), .B0(n1184), .Y(n1136) );
  INVX1 U919 ( .A(n1136), .Y(n285) );
  OA21XL U920 ( .A0(n226), .A1(n269), .B0(n1185), .Y(n1137) );
  INVX1 U921 ( .A(n1137), .Y(n270) );
  OA21XL U922 ( .A0(n174), .A1(n204), .B0(n1187), .Y(n1138) );
  INVX1 U923 ( .A(n1138), .Y(n205) );
  OA21XL U924 ( .A0(n1330), .A1(n284), .B0(n1184), .Y(n1139) );
  INVX1 U925 ( .A(n1139), .Y(n244) );
  OA21XL U926 ( .A0(n180), .A1(n204), .B0(n1186), .Y(n1140) );
  INVX1 U927 ( .A(n1140), .Y(n209) );
  OA21XL U928 ( .A0(n1328), .A1(n255), .B0(n1185), .Y(n1141) );
  INVX1 U929 ( .A(n1141), .Y(n260) );
  OA21XL U930 ( .A0(n164), .A1(n204), .B0(n1186), .Y(n1142) );
  INVX1 U931 ( .A(n1142), .Y(n216) );
  OA21XL U932 ( .A0(n223), .A1(n255), .B0(n1185), .Y(n1143) );
  INVX1 U933 ( .A(n1143), .Y(n249) );
  OA21XL U934 ( .A0(n223), .A1(n279), .B0(n1184), .Y(n1144) );
  INVX1 U935 ( .A(n1144), .Y(n277) );
  OA21XL U936 ( .A0(n155), .A1(n204), .B0(n1186), .Y(n1145) );
  INVX1 U937 ( .A(n1145), .Y(n211) );
  OA21XL U938 ( .A0(n223), .A1(n284), .B0(n1184), .Y(n1146) );
  INVX1 U939 ( .A(n1146), .Y(n282) );
  OA21XL U940 ( .A0(n223), .A1(n269), .B0(n1185), .Y(n1147) );
  INVX1 U941 ( .A(n1147), .Y(n267) );
  OA21XL U942 ( .A0(n171), .A1(n204), .B0(n1187), .Y(n1148) );
  INVX1 U943 ( .A(n1148), .Y(n202) );
  OA21XL U944 ( .A0(n1328), .A1(n284), .B0(n1184), .Y(n1149) );
  INVX1 U945 ( .A(n1149), .Y(n288) );
  OA21XL U946 ( .A0(n177), .A1(n204), .B0(n1186), .Y(n1150) );
  INVX1 U947 ( .A(n1150), .Y(n207) );
  OAI21XL U948 ( .A0(n1101), .A1(n121), .B0(n127), .Y(n1081) );
  OAI21XL U949 ( .A0(n128), .A1(n124), .B0(n121), .Y(n127) );
  OAI21XL U950 ( .A0(n1096), .A1(n121), .B0(n123), .Y(n1082) );
  OAI21XL U951 ( .A0(n124), .A1(n125), .B0(n121), .Y(n123) );
  BUFX2 U952 ( .A(n22), .Y(n1216) );
  BUFX2 U953 ( .A(n21), .Y(n1219) );
  BUFX2 U954 ( .A(n150), .Y(n1201) );
  BUFX2 U955 ( .A(n150), .Y(n1203) );
  BUFX2 U956 ( .A(n150), .Y(n1202) );
  BUFX2 U957 ( .A(n151), .Y(n1198) );
  BUFX2 U958 ( .A(n151), .Y(n1200) );
  BUFX2 U959 ( .A(n151), .Y(n1199) );
  BUFX2 U960 ( .A(n152), .Y(n1195) );
  BUFX2 U961 ( .A(n152), .Y(n1197) );
  BUFX2 U962 ( .A(n152), .Y(n1196) );
  BUFX2 U963 ( .A(n153), .Y(n1192) );
  BUFX2 U964 ( .A(n153), .Y(n1194) );
  BUFX2 U965 ( .A(n153), .Y(n1193) );
  BUFX2 U966 ( .A(n145), .Y(n1210) );
  BUFX2 U967 ( .A(n145), .Y(n1212) );
  BUFX2 U968 ( .A(n145), .Y(n1211) );
  BUFX2 U969 ( .A(n146), .Y(n1207) );
  BUFX2 U970 ( .A(n146), .Y(n1209) );
  BUFX2 U971 ( .A(n146), .Y(n1208) );
  BUFX2 U972 ( .A(n147), .Y(n1204) );
  BUFX2 U973 ( .A(n147), .Y(n1206) );
  BUFX2 U974 ( .A(n147), .Y(n1205) );
  BUFX2 U975 ( .A(n142), .Y(n1213) );
  BUFX2 U976 ( .A(n142), .Y(n1215) );
  BUFX2 U977 ( .A(n142), .Y(n1214) );
  AND2X2 U978 ( .A(n291), .B(cnt_32[2]), .Y(n266) );
  NAND2X1 U979 ( .A(n129), .B(n130), .Y(n124) );
  INVX1 U980 ( .A(n232), .Y(n1325) );
  BUFX2 U981 ( .A(n21), .Y(n1220) );
  INVX1 U982 ( .A(n1155), .Y(n1173) );
  INVX1 U983 ( .A(n1155), .Y(n1172) );
  INVX1 U984 ( .A(n1156), .Y(n1171) );
  INVX1 U985 ( .A(n1156), .Y(n1170) );
  INVX1 U986 ( .A(n1157), .Y(n1169) );
  INVX1 U987 ( .A(n1157), .Y(n1168) );
  INVX1 U988 ( .A(n1158), .Y(n1167) );
  INVX1 U989 ( .A(n1158), .Y(n1166) );
  INVX1 U990 ( .A(n1159), .Y(n1180) );
  INVX1 U991 ( .A(n1159), .Y(n1179) );
  INVX1 U992 ( .A(n1160), .Y(n1178) );
  INVX1 U993 ( .A(n1160), .Y(n1177) );
  INVX1 U994 ( .A(n1162), .Y(n1164) );
  INVX1 U995 ( .A(n1161), .Y(n1176) );
  INVX1 U996 ( .A(n1161), .Y(n1175) );
  INVX1 U997 ( .A(n1162), .Y(n1165) );
  INVX1 U998 ( .A(n226), .Y(n1327) );
  INVX1 U999 ( .A(n223), .Y(n1329) );
  BUFX2 U1000 ( .A(n29), .Y(n1163) );
  BUFX2 U1001 ( .A(n26), .Y(n1174) );
  OA21XL U1002 ( .A0(n232), .A1(n130), .B0(n1188), .Y(n132) );
  AND2X2 U1003 ( .A(n237), .B(n235), .Y(n236) );
  AO22X1 U1004 ( .A0(n1183), .A1(N94), .B0(n125), .B1(N108), .Y(n237) );
  INVX1 U1005 ( .A(n138), .Y(n1324) );
  BUFX2 U1006 ( .A(n22), .Y(n1217) );
  BUFX2 U1007 ( .A(n21), .Y(n1221) );
  BUFX2 U1008 ( .A(reset), .Y(n1271) );
  BUFX2 U1009 ( .A(clock), .Y(n1316) );
  BUFX2 U1010 ( .A(reset), .Y(n1270) );
  BUFX2 U1011 ( .A(clock), .Y(n1315) );
  BUFX2 U1012 ( .A(reset), .Y(n1269) );
  BUFX2 U1013 ( .A(clock), .Y(n1314) );
  BUFX2 U1014 ( .A(reset), .Y(n1268) );
  BUFX2 U1015 ( .A(clock), .Y(n1313) );
  BUFX2 U1016 ( .A(reset), .Y(n1272) );
  AND4X1 U1017 ( .A(n8), .B(n9), .C(n10), .D(n11), .Y(n734) );
  AOI222XL U1018 ( .A0(n1321), .A1(n1091), .B0(n1327), .B1(n15), .C0(n1329), 
        .C1(n17), .Y(n11) );
  OAI21XL U1019 ( .A0(n24), .A1(n25), .B0(n1174), .Y(n10) );
  OAI21XL U1020 ( .A0(n27), .A1(n28), .B0(n1163), .Y(n8) );
  AND4X1 U1021 ( .A(n30), .B(n9), .C(n31), .D(n32), .Y(n783) );
  AOI222XL U1022 ( .A0(n1321), .A1(n1092), .B0(n1327), .B1(n34), .C0(n1329), 
        .C1(n35), .Y(n32) );
  OAI21XL U1023 ( .A0(n38), .A1(n39), .B0(n1174), .Y(n31) );
  OAI21XL U1024 ( .A0(n40), .A1(n41), .B0(n1163), .Y(n30) );
  AND4X1 U1025 ( .A(n42), .B(n9), .C(n43), .D(n44), .Y(n832) );
  AOI222XL U1026 ( .A0(n1181), .A1(n1093), .B0(n1327), .B1(n46), .C0(n1329), 
        .C1(n47), .Y(n44) );
  OAI21XL U1027 ( .A0(n50), .A1(n51), .B0(n1174), .Y(n43) );
  OAI21XL U1028 ( .A0(n52), .A1(n53), .B0(n1163), .Y(n42) );
  AND4X1 U1029 ( .A(n54), .B(n9), .C(n55), .D(n56), .Y(n881) );
  AOI222XL U1030 ( .A0(n1321), .A1(n1095), .B0(n1327), .B1(n58), .C0(n1329), 
        .C1(n59), .Y(n56) );
  OAI21XL U1031 ( .A0(n62), .A1(n63), .B0(n1174), .Y(n55) );
  OAI21XL U1032 ( .A0(n64), .A1(n65), .B0(n1163), .Y(n54) );
  AND4X1 U1033 ( .A(n66), .B(n9), .C(n67), .D(n68), .Y(n930) );
  AOI222XL U1034 ( .A0(n1181), .A1(n1094), .B0(n1327), .B1(n70), .C0(n1329), 
        .C1(n71), .Y(n68) );
  OAI21XL U1035 ( .A0(n74), .A1(n75), .B0(n1174), .Y(n67) );
  OAI21XL U1036 ( .A0(n76), .A1(n77), .B0(n1163), .Y(n66) );
  AND4X1 U1037 ( .A(n78), .B(n9), .C(n79), .D(n80), .Y(n979) );
  AOI222XL U1038 ( .A0(n1321), .A1(n1100), .B0(n1327), .B1(n82), .C0(n1329), 
        .C1(n83), .Y(n80) );
  OAI21XL U1039 ( .A0(n86), .A1(n87), .B0(n1174), .Y(n79) );
  OAI21XL U1040 ( .A0(n88), .A1(n89), .B0(n1163), .Y(n78) );
  AND4X1 U1041 ( .A(n102), .B(n9), .C(n103), .D(n104), .Y(n1028) );
  AOI222XL U1042 ( .A0(n1181), .A1(n1098), .B0(n1327), .B1(n106), .C0(n1329), 
        .C1(n107), .Y(n104) );
  OAI21XL U1043 ( .A0(n110), .A1(n111), .B0(n1174), .Y(n103) );
  OAI21XL U1044 ( .A0(n114), .A1(n115), .B0(n1163), .Y(n102) );
  AND4X1 U1045 ( .A(n90), .B(n9), .C(n91), .D(n92), .Y(n1087) );
  AOI222XL U1046 ( .A0(n1321), .A1(n1099), .B0(n1327), .B1(n94), .C0(n1329), 
        .C1(n95), .Y(n92) );
  OAI21XL U1047 ( .A0(n98), .A1(n99), .B0(n1174), .Y(n91) );
  OAI21XL U1048 ( .A0(n100), .A1(n101), .B0(n1163), .Y(n90) );
  BUFX2 U1049 ( .A(n22), .Y(n1218) );
  OAI2BB2XL U1050 ( .B0(n1191), .B1(n1095), .A0N(data[4]), .A1N(n1089), .Y(
        display_data[4]) );
  INVX1 U1051 ( .A(data[0]), .Y(n1332) );
  INVX1 U1052 ( .A(data[1]), .Y(n1326) );
  OR2X1 U1053 ( .A(ready), .B(result_valid), .Y(_8_net_) );
  NAND2X1 U1054 ( .A(n128), .B(phase[0]), .Y(n129) );
  NOR2X1 U1055 ( .A(phase[1]), .B(phase[2]), .Y(n128) );
  NOR4X1 U1056 ( .A(next_status[2]), .B(next_status[0]), .C(n1096), .D(n239), 
        .Y(N58) );
  NOR4X1 U1057 ( .A(next_status[2]), .B(n1101), .C(n1096), .D(n129), .Y(N57)
         );
  NOR2BX1 U1058 ( .AN(phase[1]), .B(phase[0]), .Y(n233) );
  OR3X2 U1059 ( .A(n1151), .B(n1152), .C(n1153), .Y(n232) );
  XOR2X1 U1060 ( .A(next_status[2]), .B(phase[2]), .Y(n1151) );
  XOR2X1 U1061 ( .A(next_status[0]), .B(phase[0]), .Y(n1152) );
  XOR2X1 U1062 ( .A(next_status[1]), .B(phase[1]), .Y(n1153) );
  NAND3BX1 U1063 ( .AN(phase[0]), .B(n128), .C(n1325), .Y(n138) );
  OAI22XL U1064 ( .A0(result[39]), .A1(n1223), .B0(result[7]), .B1(n1226), .Y(
        n27) );
  OAI22XL U1065 ( .A0(result[47]), .A1(n1223), .B0(result[15]), .B1(n1226), 
        .Y(n24) );
  OAI22XL U1066 ( .A0(result[38]), .A1(n1223), .B0(result[6]), .B1(n1226), .Y(
        n40) );
  OAI22XL U1067 ( .A0(result[46]), .A1(n1223), .B0(result[14]), .B1(n1226), 
        .Y(n38) );
  OAI22XL U1068 ( .A0(result[37]), .A1(n1222), .B0(result[5]), .B1(n1225), .Y(
        n52) );
  OAI22XL U1069 ( .A0(result[45]), .A1(n1223), .B0(result[13]), .B1(n1226), 
        .Y(n50) );
  OAI22XL U1070 ( .A0(result[36]), .A1(n1223), .B0(result[4]), .B1(n1226), .Y(
        n64) );
  OAI22XL U1071 ( .A0(result[44]), .A1(n1222), .B0(result[12]), .B1(n1225), 
        .Y(n62) );
  OAI22XL U1072 ( .A0(result[35]), .A1(n1222), .B0(result[3]), .B1(n1225), .Y(
        n76) );
  OAI22XL U1073 ( .A0(result[43]), .A1(n1222), .B0(result[11]), .B1(n1225), 
        .Y(n74) );
  OAI22XL U1074 ( .A0(result[34]), .A1(n1222), .B0(result[2]), .B1(n1225), .Y(
        n88) );
  OAI22XL U1075 ( .A0(result[42]), .A1(n1222), .B0(result[10]), .B1(n1225), 
        .Y(n86) );
  OAI22XL U1076 ( .A0(result[32]), .A1(n1222), .B0(result[0]), .B1(n1225), .Y(
        n114) );
  OAI22XL U1077 ( .A0(result[40]), .A1(n1222), .B0(result[8]), .B1(n1225), .Y(
        n110) );
  OAI22XL U1078 ( .A0(result[33]), .A1(n1222), .B0(result[1]), .B1(n1225), .Y(
        n100) );
  OAI22XL U1079 ( .A0(result[41]), .A1(n1222), .B0(result[9]), .B1(n1225), .Y(
        n98) );
  OAI22XL U1080 ( .A0(result[103]), .A1(n1218), .B0(result[71]), .B1(n1220), 
        .Y(n28) );
  OAI22XL U1081 ( .A0(result[111]), .A1(n1218), .B0(result[79]), .B1(n1220), 
        .Y(n25) );
  OAI22XL U1082 ( .A0(result[102]), .A1(n22), .B0(result[70]), .B1(n1220), .Y(
        n41) );
  OAI22XL U1083 ( .A0(result[110]), .A1(n1218), .B0(result[78]), .B1(n1220), 
        .Y(n39) );
  OAI22XL U1084 ( .A0(result[101]), .A1(n1216), .B0(result[69]), .B1(n1219), 
        .Y(n53) );
  OAI22XL U1085 ( .A0(result[109]), .A1(n22), .B0(result[77]), .B1(n1220), .Y(
        n51) );
  OAI22XL U1086 ( .A0(result[100]), .A1(n1218), .B0(result[68]), .B1(n1220), 
        .Y(n65) );
  OAI22XL U1087 ( .A0(result[108]), .A1(n1216), .B0(result[76]), .B1(n1219), 
        .Y(n63) );
  OAI22XL U1088 ( .A0(result[99]), .A1(n1216), .B0(result[67]), .B1(n1219), 
        .Y(n77) );
  OAI22XL U1089 ( .A0(result[107]), .A1(n1216), .B0(result[75]), .B1(n1219), 
        .Y(n75) );
  OAI22XL U1090 ( .A0(result[98]), .A1(n1216), .B0(result[66]), .B1(n1219), 
        .Y(n89) );
  OAI22XL U1091 ( .A0(result[106]), .A1(n1216), .B0(result[74]), .B1(n1219), 
        .Y(n87) );
  OAI22XL U1092 ( .A0(result[96]), .A1(n1216), .B0(result[64]), .B1(n1219), 
        .Y(n115) );
  OAI22XL U1093 ( .A0(result[104]), .A1(n1216), .B0(result[72]), .B1(n1219), 
        .Y(n111) );
  OAI22XL U1094 ( .A0(result[97]), .A1(n1216), .B0(result[65]), .B1(n1219), 
        .Y(n101) );
  OAI22XL U1095 ( .A0(result[105]), .A1(n1216), .B0(result[73]), .B1(n1219), 
        .Y(n99) );
  NAND2X1 U1096 ( .A(n683), .B(n117), .Y(n22) );
  NAND2X1 U1097 ( .A(n683), .B(n116), .Y(n21) );
  OAI22XL U1098 ( .A0(n295), .A1(n186), .B0(n1125), .B1(n1202), .Y(n686) );
  OAI22XL U1099 ( .A0(n296), .A1(n192), .B0(n1126), .B1(n1202), .Y(n687) );
  OAI22XL U1100 ( .A0(n297), .A1(n196), .B0(n1124), .B1(n1202), .Y(n688) );
  OAI22XL U1101 ( .A0(n298), .A1(n200), .B0(n1123), .B1(n1202), .Y(n689) );
  OAI22XL U1102 ( .A0(n299), .A1(n205), .B0(n1138), .B1(n1203), .Y(n690) );
  OAI22XL U1103 ( .A0(n300), .A1(n209), .B0(n1140), .B1(n1203), .Y(n691) );
  OAI22XL U1104 ( .A0(n301), .A1(n214), .B0(n1135), .B1(n1203), .Y(n692) );
  OAI22XL U1105 ( .A0(n302), .A1(n218), .B0(n1132), .B1(n1203), .Y(n693) );
  OAI22XL U1106 ( .A0(n303), .A1(n224), .B0(n1117), .B1(n1203), .Y(n694) );
  OAI22XL U1107 ( .A0(n304), .A1(n143), .B0(n1121), .B1(n150), .Y(n695) );
  OAI22XL U1108 ( .A0(n305), .A1(n157), .B0(n1116), .B1(n1201), .Y(n696) );
  OAI22XL U1109 ( .A0(n306), .A1(n165), .B0(n1115), .B1(n1201), .Y(n697) );
  OAI22XL U1110 ( .A0(n307), .A1(n172), .B0(n1105), .B1(n1201), .Y(n698) );
  OAI22XL U1111 ( .A0(n308), .A1(n178), .B0(n1106), .B1(n1201), .Y(n699) );
  OAI22XL U1112 ( .A0(n309), .A1(n188), .B0(n1104), .B1(n1202), .Y(n700) );
  OAI22XL U1113 ( .A0(n310), .A1(n160), .B0(n1103), .B1(n1201), .Y(n701) );
  OAI22XL U1114 ( .A0(n311), .A1(n140), .B0(n1107), .B1(n1203), .Y(n702) );
  OAI22XL U1115 ( .A0(n312), .A1(n181), .B0(n1108), .B1(n1201), .Y(n703) );
  OAI22XL U1116 ( .A0(n313), .A1(n175), .B0(n1113), .B1(n1201), .Y(n704) );
  OAI22XL U1117 ( .A0(n314), .A1(n168), .B0(n1111), .B1(n1201), .Y(n705) );
  OAI22XL U1118 ( .A0(n315), .A1(n162), .B0(n1122), .B1(n1201), .Y(n706) );
  OAI22XL U1119 ( .A0(n316), .A1(n148), .B0(n1118), .B1(n1201), .Y(n707) );
  OAI22XL U1120 ( .A0(n317), .A1(n227), .B0(n1120), .B1(n150), .Y(n708) );
  OAI22XL U1121 ( .A0(n318), .A1(n220), .B0(n1119), .B1(n1203), .Y(n709) );
  OAI22XL U1122 ( .A0(n319), .A1(n216), .B0(n1142), .B1(n1203), .Y(n710) );
  OAI22XL U1123 ( .A0(n320), .A1(n211), .B0(n1145), .B1(n1203), .Y(n711) );
  OAI22XL U1124 ( .A0(n321), .A1(n207), .B0(n1150), .B1(n1203), .Y(n712) );
  OAI22XL U1125 ( .A0(n322), .A1(n202), .B0(n1148), .B1(n1202), .Y(n713) );
  OAI22XL U1126 ( .A0(n323), .A1(n198), .B0(n1127), .B1(n1202), .Y(n714) );
  OAI22XL U1127 ( .A0(n324), .A1(n194), .B0(n1128), .B1(n1202), .Y(n715) );
  OAI22XL U1128 ( .A0(n325), .A1(n190), .B0(n1130), .B1(n1202), .Y(n716) );
  OAI22XL U1129 ( .A0(n326), .A1(n183), .B0(n1129), .B1(n1202), .Y(n717) );
  OAI22XL U1130 ( .A0(n327), .A1(n285), .B0(n1136), .B1(n1173), .Y(n718) );
  OAI22XL U1131 ( .A0(n328), .A1(n244), .B0(n1139), .B1(n1173), .Y(n719) );
  OAI22XL U1132 ( .A0(n329), .A1(n256), .B0(n1133), .B1(n1173), .Y(n720) );
  OAI22XL U1133 ( .A0(n330), .A1(n263), .B0(n1131), .B1(n1172), .Y(n721) );
  OAI22XL U1134 ( .A0(n331), .A1(n270), .B0(n1137), .B1(n1172), .Y(n722) );
  OAI22XL U1135 ( .A0(n332), .A1(n274), .B0(n1109), .B1(n1172), .Y(n723) );
  OAI22XL U1136 ( .A0(n333), .A1(n280), .B0(n1134), .B1(n1172), .Y(n724) );
  OAI22XL U1137 ( .A0(n334), .A1(n258), .B0(n1114), .B1(n1172), .Y(n725) );
  OAI22XL U1138 ( .A0(n335), .A1(n241), .B0(n1110), .B1(n1173), .Y(n726) );
  OAI22XL U1139 ( .A0(n336), .A1(n277), .B0(n1144), .B1(n1173), .Y(n727) );
  OAI22XL U1140 ( .A0(n337), .A1(n272), .B0(n1112), .B1(n1173), .Y(n728) );
  OAI22XL U1141 ( .A0(n338), .A1(n267), .B0(n1147), .B1(n1173), .Y(n729) );
  OAI22XL U1142 ( .A0(n339), .A1(n260), .B0(n1141), .B1(n1173), .Y(n730) );
  OAI22XL U1143 ( .A0(n340), .A1(n249), .B0(n1143), .B1(n1172), .Y(n731) );
  OAI22XL U1144 ( .A0(n341), .A1(n288), .B0(n1149), .B1(n1172), .Y(n732) );
  OAI22XL U1145 ( .A0(n342), .A1(n282), .B0(n1146), .B1(n1172), .Y(n733) );
  OAI22XL U1146 ( .A0(n343), .A1(n186), .B0(n1125), .B1(n1199), .Y(n735) );
  OAI22XL U1147 ( .A0(n344), .A1(n192), .B0(n1126), .B1(n1199), .Y(n736) );
  OAI22XL U1148 ( .A0(n345), .A1(n196), .B0(n1124), .B1(n1199), .Y(n737) );
  OAI22XL U1149 ( .A0(n346), .A1(n200), .B0(n1123), .B1(n1199), .Y(n738) );
  OAI22XL U1150 ( .A0(n347), .A1(n205), .B0(n1138), .B1(n1200), .Y(n739) );
  OAI22XL U1151 ( .A0(n348), .A1(n209), .B0(n1140), .B1(n1200), .Y(n740) );
  OAI22XL U1152 ( .A0(n349), .A1(n214), .B0(n1135), .B1(n1200), .Y(n741) );
  OAI22XL U1153 ( .A0(n350), .A1(n218), .B0(n1132), .B1(n1200), .Y(n742) );
  OAI22XL U1154 ( .A0(n351), .A1(n224), .B0(n1117), .B1(n1200), .Y(n743) );
  OAI22XL U1155 ( .A0(n352), .A1(n143), .B0(n1121), .B1(n151), .Y(n744) );
  OAI22XL U1156 ( .A0(n353), .A1(n157), .B0(n1116), .B1(n1198), .Y(n745) );
  OAI22XL U1157 ( .A0(n354), .A1(n165), .B0(n1115), .B1(n1198), .Y(n746) );
  OAI22XL U1158 ( .A0(n356), .A1(n178), .B0(n1106), .B1(n1198), .Y(n748) );
  OAI22XL U1159 ( .A0(n357), .A1(n188), .B0(n1104), .B1(n1199), .Y(n749) );
  OAI22XL U1160 ( .A0(n358), .A1(n160), .B0(n1103), .B1(n1198), .Y(n750) );
  OAI22XL U1161 ( .A0(n359), .A1(n140), .B0(n1107), .B1(n1200), .Y(n751) );
  OAI22XL U1162 ( .A0(n360), .A1(n181), .B0(n1108), .B1(n1198), .Y(n752) );
  OAI22XL U1163 ( .A0(n361), .A1(n175), .B0(n1113), .B1(n1198), .Y(n753) );
  OAI22XL U1164 ( .A0(n362), .A1(n168), .B0(n1111), .B1(n1198), .Y(n754) );
  OAI22XL U1165 ( .A0(n364), .A1(n148), .B0(n1118), .B1(n1198), .Y(n756) );
  OAI22XL U1166 ( .A0(n365), .A1(n227), .B0(n1120), .B1(n151), .Y(n757) );
  OAI22XL U1167 ( .A0(n366), .A1(n220), .B0(n1119), .B1(n1200), .Y(n758) );
  OAI22XL U1168 ( .A0(n367), .A1(n216), .B0(n1142), .B1(n1200), .Y(n759) );
  OAI22XL U1169 ( .A0(n368), .A1(n211), .B0(n1145), .B1(n1200), .Y(n760) );
  OAI22XL U1170 ( .A0(n369), .A1(n207), .B0(n1150), .B1(n1200), .Y(n761) );
  OAI22XL U1171 ( .A0(n370), .A1(n202), .B0(n1148), .B1(n1199), .Y(n762) );
  OAI22XL U1172 ( .A0(n371), .A1(n198), .B0(n1127), .B1(n1199), .Y(n763) );
  OAI22XL U1173 ( .A0(n372), .A1(n194), .B0(n1128), .B1(n1199), .Y(n764) );
  OAI22XL U1174 ( .A0(n373), .A1(n190), .B0(n1130), .B1(n1199), .Y(n765) );
  OAI22XL U1175 ( .A0(n374), .A1(n183), .B0(n1129), .B1(n1199), .Y(n766) );
  OAI22XL U1176 ( .A0(n375), .A1(n285), .B0(n1136), .B1(n1171), .Y(n767) );
  OAI22XL U1177 ( .A0(n376), .A1(n244), .B0(n1139), .B1(n1171), .Y(n768) );
  OAI22XL U1178 ( .A0(n377), .A1(n256), .B0(n1133), .B1(n1171), .Y(n769) );
  OAI22XL U1179 ( .A0(n378), .A1(n263), .B0(n1131), .B1(n1171), .Y(n770) );
  OAI22XL U1180 ( .A0(n379), .A1(n270), .B0(n1137), .B1(n1170), .Y(n771) );
  OAI22XL U1181 ( .A0(n380), .A1(n274), .B0(n1109), .B1(n1170), .Y(n772) );
  OAI22XL U1182 ( .A0(n381), .A1(n280), .B0(n1134), .B1(n1170), .Y(n773) );
  OAI22XL U1183 ( .A0(n382), .A1(n258), .B0(n1114), .B1(n1170), .Y(n774) );
  OAI22XL U1184 ( .A0(n383), .A1(n241), .B0(n1110), .B1(n1171), .Y(n775) );
  OAI22XL U1185 ( .A0(n384), .A1(n277), .B0(n1144), .B1(n1171), .Y(n776) );
  OAI22XL U1186 ( .A0(n385), .A1(n272), .B0(n1112), .B1(n1171), .Y(n777) );
  OAI22XL U1187 ( .A0(n386), .A1(n267), .B0(n1147), .B1(n1171), .Y(n778) );
  OAI22XL U1188 ( .A0(n387), .A1(n260), .B0(n1141), .B1(n1170), .Y(n779) );
  OAI22XL U1189 ( .A0(n388), .A1(n249), .B0(n1143), .B1(n1170), .Y(n780) );
  OAI22XL U1190 ( .A0(n389), .A1(n288), .B0(n1149), .B1(n1170), .Y(n781) );
  OAI22XL U1191 ( .A0(n390), .A1(n282), .B0(n1146), .B1(n1170), .Y(n782) );
  OAI22XL U1192 ( .A0(n391), .A1(n186), .B0(n1125), .B1(n1196), .Y(n784) );
  OAI22XL U1193 ( .A0(n392), .A1(n192), .B0(n1126), .B1(n1196), .Y(n785) );
  OAI22XL U1194 ( .A0(n393), .A1(n196), .B0(n1124), .B1(n1196), .Y(n786) );
  OAI22XL U1195 ( .A0(n394), .A1(n200), .B0(n1123), .B1(n1196), .Y(n787) );
  OAI22XL U1196 ( .A0(n395), .A1(n205), .B0(n1138), .B1(n1197), .Y(n788) );
  OAI22XL U1197 ( .A0(n396), .A1(n209), .B0(n1140), .B1(n1197), .Y(n789) );
  OAI22XL U1198 ( .A0(n397), .A1(n214), .B0(n1135), .B1(n1197), .Y(n790) );
  OAI22XL U1199 ( .A0(n398), .A1(n218), .B0(n1132), .B1(n1197), .Y(n791) );
  OAI22XL U1200 ( .A0(n399), .A1(n224), .B0(n1117), .B1(n1197), .Y(n792) );
  OAI22XL U1201 ( .A0(n400), .A1(n143), .B0(n1121), .B1(n152), .Y(n793) );
  OAI22XL U1202 ( .A0(n401), .A1(n157), .B0(n1116), .B1(n1195), .Y(n794) );
  OAI22XL U1203 ( .A0(n402), .A1(n165), .B0(n1115), .B1(n1195), .Y(n795) );
  OAI22XL U1204 ( .A0(n403), .A1(n172), .B0(n1105), .B1(n1195), .Y(n796) );
  OAI22XL U1205 ( .A0(n404), .A1(n178), .B0(n1106), .B1(n1195), .Y(n797) );
  OAI22XL U1206 ( .A0(n405), .A1(n188), .B0(n1104), .B1(n1196), .Y(n798) );
  OAI22XL U1207 ( .A0(n406), .A1(n160), .B0(n1103), .B1(n1195), .Y(n799) );
  OAI22XL U1208 ( .A0(n407), .A1(n140), .B0(n1107), .B1(n1197), .Y(n800) );
  OAI22XL U1209 ( .A0(n408), .A1(n181), .B0(n1108), .B1(n1195), .Y(n801) );
  OAI22XL U1210 ( .A0(n409), .A1(n175), .B0(n1113), .B1(n1195), .Y(n802) );
  OAI22XL U1211 ( .A0(n410), .A1(n168), .B0(n1111), .B1(n1195), .Y(n803) );
  OAI22XL U1212 ( .A0(n411), .A1(n162), .B0(n1122), .B1(n1195), .Y(n804) );
  OAI22XL U1213 ( .A0(n412), .A1(n148), .B0(n1118), .B1(n1195), .Y(n805) );
  OAI22XL U1214 ( .A0(n413), .A1(n227), .B0(n1120), .B1(n152), .Y(n806) );
  OAI22XL U1215 ( .A0(n414), .A1(n220), .B0(n1119), .B1(n1197), .Y(n807) );
  OAI22XL U1216 ( .A0(n415), .A1(n216), .B0(n1142), .B1(n1197), .Y(n808) );
  OAI22XL U1217 ( .A0(n416), .A1(n211), .B0(n1145), .B1(n1197), .Y(n809) );
  OAI22XL U1218 ( .A0(n417), .A1(n207), .B0(n1150), .B1(n1197), .Y(n810) );
  OAI22XL U1219 ( .A0(n418), .A1(n202), .B0(n1148), .B1(n1196), .Y(n811) );
  OAI22XL U1220 ( .A0(n419), .A1(n198), .B0(n1127), .B1(n1196), .Y(n812) );
  OAI22XL U1221 ( .A0(n420), .A1(n194), .B0(n1128), .B1(n1196), .Y(n813) );
  OAI22XL U1222 ( .A0(n421), .A1(n190), .B0(n1130), .B1(n1196), .Y(n814) );
  OAI22XL U1223 ( .A0(n422), .A1(n183), .B0(n1129), .B1(n1196), .Y(n815) );
  OAI22XL U1224 ( .A0(n423), .A1(n285), .B0(n1136), .B1(n1169), .Y(n816) );
  OAI22XL U1225 ( .A0(n424), .A1(n244), .B0(n1139), .B1(n1169), .Y(n817) );
  OAI22XL U1226 ( .A0(n425), .A1(n256), .B0(n1133), .B1(n1169), .Y(n818) );
  OAI22XL U1227 ( .A0(n426), .A1(n263), .B0(n1131), .B1(n1169), .Y(n819) );
  OAI22XL U1228 ( .A0(n427), .A1(n270), .B0(n1137), .B1(n1168), .Y(n820) );
  OAI22XL U1229 ( .A0(n428), .A1(n274), .B0(n1109), .B1(n1168), .Y(n821) );
  OAI22XL U1230 ( .A0(n429), .A1(n280), .B0(n1134), .B1(n1168), .Y(n822) );
  OAI22XL U1231 ( .A0(n430), .A1(n258), .B0(n1114), .B1(n1169), .Y(n823) );
  OAI22XL U1232 ( .A0(n431), .A1(n241), .B0(n1110), .B1(n1169), .Y(n824) );
  OAI22XL U1233 ( .A0(n432), .A1(n277), .B0(n1144), .B1(n1169), .Y(n825) );
  OAI22XL U1234 ( .A0(n433), .A1(n272), .B0(n1112), .B1(n1169), .Y(n826) );
  OAI22XL U1235 ( .A0(n434), .A1(n267), .B0(n1147), .B1(n1168), .Y(n827) );
  OAI22XL U1236 ( .A0(n435), .A1(n260), .B0(n1141), .B1(n1168), .Y(n828) );
  OAI22XL U1237 ( .A0(n436), .A1(n249), .B0(n1143), .B1(n1168), .Y(n829) );
  OAI22XL U1238 ( .A0(n437), .A1(n288), .B0(n1149), .B1(n1168), .Y(n830) );
  OAI22XL U1239 ( .A0(n438), .A1(n282), .B0(n1146), .B1(n1168), .Y(n831) );
  OAI22XL U1240 ( .A0(n439), .A1(n186), .B0(n1125), .B1(n1193), .Y(n833) );
  OAI22XL U1241 ( .A0(n440), .A1(n192), .B0(n1126), .B1(n1193), .Y(n834) );
  OAI22XL U1242 ( .A0(n441), .A1(n196), .B0(n1124), .B1(n1193), .Y(n835) );
  OAI22XL U1243 ( .A0(n442), .A1(n200), .B0(n1123), .B1(n1193), .Y(n836) );
  OAI22XL U1244 ( .A0(n443), .A1(n205), .B0(n1138), .B1(n1194), .Y(n837) );
  OAI22XL U1245 ( .A0(n444), .A1(n209), .B0(n1140), .B1(n1194), .Y(n838) );
  OAI22XL U1246 ( .A0(n445), .A1(n214), .B0(n1135), .B1(n1194), .Y(n839) );
  OAI22XL U1247 ( .A0(n446), .A1(n218), .B0(n1132), .B1(n1194), .Y(n840) );
  OAI22XL U1248 ( .A0(n447), .A1(n224), .B0(n1117), .B1(n1194), .Y(n841) );
  OAI22XL U1249 ( .A0(n448), .A1(n143), .B0(n1121), .B1(n153), .Y(n842) );
  OAI22XL U1250 ( .A0(n449), .A1(n157), .B0(n1116), .B1(n1192), .Y(n843) );
  OAI22XL U1251 ( .A0(n450), .A1(n165), .B0(n1115), .B1(n1192), .Y(n844) );
  OAI22XL U1252 ( .A0(n451), .A1(n172), .B0(n1105), .B1(n1192), .Y(n845) );
  OAI22XL U1253 ( .A0(n452), .A1(n178), .B0(n1106), .B1(n1192), .Y(n846) );
  OAI22XL U1254 ( .A0(n453), .A1(n188), .B0(n1104), .B1(n1193), .Y(n847) );
  OAI22XL U1255 ( .A0(n454), .A1(n160), .B0(n1103), .B1(n1192), .Y(n848) );
  OAI22XL U1256 ( .A0(n455), .A1(n140), .B0(n1107), .B1(n1194), .Y(n849) );
  OAI22XL U1257 ( .A0(n456), .A1(n181), .B0(n1108), .B1(n1192), .Y(n850) );
  OAI22XL U1258 ( .A0(n457), .A1(n175), .B0(n1113), .B1(n1192), .Y(n851) );
  OAI22XL U1259 ( .A0(n458), .A1(n168), .B0(n1111), .B1(n1192), .Y(n852) );
  OAI22XL U1260 ( .A0(n459), .A1(n162), .B0(n1122), .B1(n1192), .Y(n853) );
  OAI22XL U1261 ( .A0(n460), .A1(n148), .B0(n1118), .B1(n1192), .Y(n854) );
  OAI22XL U1262 ( .A0(n461), .A1(n227), .B0(n1120), .B1(n153), .Y(n855) );
  OAI22XL U1263 ( .A0(n462), .A1(n220), .B0(n1119), .B1(n1194), .Y(n856) );
  OAI22XL U1264 ( .A0(n463), .A1(n216), .B0(n1142), .B1(n1194), .Y(n857) );
  OAI22XL U1265 ( .A0(n464), .A1(n211), .B0(n1145), .B1(n1194), .Y(n858) );
  OAI22XL U1266 ( .A0(n465), .A1(n207), .B0(n1150), .B1(n1194), .Y(n859) );
  OAI22XL U1267 ( .A0(n466), .A1(n202), .B0(n1148), .B1(n1193), .Y(n860) );
  OAI22XL U1268 ( .A0(n467), .A1(n198), .B0(n1127), .B1(n1193), .Y(n861) );
  OAI22XL U1269 ( .A0(n468), .A1(n194), .B0(n1128), .B1(n1193), .Y(n862) );
  OAI22XL U1270 ( .A0(n469), .A1(n190), .B0(n1130), .B1(n1193), .Y(n863) );
  OAI22XL U1271 ( .A0(n470), .A1(n183), .B0(n1129), .B1(n1193), .Y(n864) );
  OAI22XL U1272 ( .A0(n471), .A1(n285), .B0(n1136), .B1(n1167), .Y(n865) );
  OAI22XL U1273 ( .A0(n472), .A1(n244), .B0(n1139), .B1(n1167), .Y(n866) );
  OAI22XL U1274 ( .A0(n473), .A1(n256), .B0(n1133), .B1(n1167), .Y(n867) );
  OAI22XL U1275 ( .A0(n474), .A1(n263), .B0(n1131), .B1(n1167), .Y(n868) );
  OAI22XL U1276 ( .A0(n475), .A1(n270), .B0(n1137), .B1(n1167), .Y(n869) );
  OAI22XL U1277 ( .A0(n476), .A1(n274), .B0(n1109), .B1(n1166), .Y(n870) );
  OAI22XL U1278 ( .A0(n477), .A1(n280), .B0(n1134), .B1(n1166), .Y(n871) );
  OAI22XL U1279 ( .A0(n478), .A1(n258), .B0(n1114), .B1(n1166), .Y(n872) );
  OAI22XL U1280 ( .A0(n479), .A1(n241), .B0(n1110), .B1(n1167), .Y(n873) );
  OAI22XL U1281 ( .A0(n480), .A1(n277), .B0(n1144), .B1(n1167), .Y(n874) );
  OAI22XL U1282 ( .A0(n481), .A1(n272), .B0(n1112), .B1(n1167), .Y(n875) );
  OAI22XL U1283 ( .A0(n482), .A1(n267), .B0(n1147), .B1(n1166), .Y(n876) );
  OAI22XL U1284 ( .A0(n483), .A1(n260), .B0(n1141), .B1(n1166), .Y(n877) );
  OAI22XL U1285 ( .A0(n484), .A1(n249), .B0(n1143), .B1(n1166), .Y(n878) );
  OAI22XL U1286 ( .A0(n485), .A1(n288), .B0(n1149), .B1(n1166), .Y(n879) );
  OAI22XL U1287 ( .A0(n486), .A1(n282), .B0(n1146), .B1(n1166), .Y(n880) );
  OAI22XL U1288 ( .A0(n487), .A1(n186), .B0(n1125), .B1(n1211), .Y(n882) );
  OAI22XL U1289 ( .A0(n488), .A1(n192), .B0(n1126), .B1(n1211), .Y(n883) );
  OAI22XL U1290 ( .A0(n489), .A1(n196), .B0(n1124), .B1(n1211), .Y(n884) );
  OAI22XL U1291 ( .A0(n490), .A1(n200), .B0(n1123), .B1(n1211), .Y(n885) );
  OAI22XL U1292 ( .A0(n491), .A1(n205), .B0(n1138), .B1(n1212), .Y(n886) );
  OAI22XL U1293 ( .A0(n492), .A1(n209), .B0(n1140), .B1(n1212), .Y(n887) );
  OAI22XL U1294 ( .A0(n493), .A1(n214), .B0(n1135), .B1(n1212), .Y(n888) );
  OAI22XL U1295 ( .A0(n494), .A1(n218), .B0(n1132), .B1(n1212), .Y(n889) );
  OAI22XL U1296 ( .A0(n495), .A1(n224), .B0(n1117), .B1(n145), .Y(n890) );
  OAI22XL U1297 ( .A0(n496), .A1(n143), .B0(n1121), .B1(n1210), .Y(n891) );
  OAI22XL U1298 ( .A0(n497), .A1(n157), .B0(n1116), .B1(n1210), .Y(n892) );
  OAI22XL U1299 ( .A0(n498), .A1(n165), .B0(n1115), .B1(n1210), .Y(n893) );
  OAI22XL U1300 ( .A0(n499), .A1(n172), .B0(n1105), .B1(n1210), .Y(n894) );
  OAI22XL U1301 ( .A0(n500), .A1(n178), .B0(n1106), .B1(n1210), .Y(n895) );
  OAI22XL U1302 ( .A0(n501), .A1(n188), .B0(n1104), .B1(n1211), .Y(n896) );
  OAI22XL U1303 ( .A0(n502), .A1(n160), .B0(n1103), .B1(n1210), .Y(n897) );
  OAI22XL U1304 ( .A0(n503), .A1(n140), .B0(n1107), .B1(n1212), .Y(n898) );
  OAI22XL U1305 ( .A0(n504), .A1(n181), .B0(n1108), .B1(n1211), .Y(n899) );
  OAI22XL U1306 ( .A0(n505), .A1(n175), .B0(n1113), .B1(n1210), .Y(n900) );
  OAI22XL U1307 ( .A0(n506), .A1(n168), .B0(n1111), .B1(n1210), .Y(n901) );
  OAI22XL U1308 ( .A0(n507), .A1(n162), .B0(n1122), .B1(n1210), .Y(n902) );
  OAI22XL U1309 ( .A0(n508), .A1(n148), .B0(n1118), .B1(n1210), .Y(n903) );
  OAI22XL U1310 ( .A0(n509), .A1(n227), .B0(n1120), .B1(n145), .Y(n904) );
  OAI22XL U1311 ( .A0(n510), .A1(n220), .B0(n1119), .B1(n1212), .Y(n905) );
  OAI22XL U1312 ( .A0(n511), .A1(n216), .B0(n1142), .B1(n1212), .Y(n906) );
  OAI22XL U1313 ( .A0(n512), .A1(n211), .B0(n1145), .B1(n1212), .Y(n907) );
  OAI22XL U1314 ( .A0(n513), .A1(n207), .B0(n1150), .B1(n1212), .Y(n908) );
  OAI22XL U1315 ( .A0(n514), .A1(n202), .B0(n1148), .B1(n1212), .Y(n909) );
  OAI22XL U1316 ( .A0(n515), .A1(n198), .B0(n1127), .B1(n1211), .Y(n910) );
  OAI22XL U1317 ( .A0(n516), .A1(n194), .B0(n1128), .B1(n1211), .Y(n911) );
  OAI22XL U1318 ( .A0(n517), .A1(n190), .B0(n1130), .B1(n1211), .Y(n912) );
  OAI22XL U1319 ( .A0(n518), .A1(n183), .B0(n1129), .B1(n1211), .Y(n913) );
  OAI22XL U1320 ( .A0(n519), .A1(n285), .B0(n1136), .B1(n1179), .Y(n914) );
  OAI22XL U1321 ( .A0(n520), .A1(n244), .B0(n1139), .B1(n1179), .Y(n915) );
  OAI22XL U1322 ( .A0(n521), .A1(n256), .B0(n1133), .B1(n1179), .Y(n916) );
  OAI22XL U1323 ( .A0(n522), .A1(n263), .B0(n1131), .B1(n1179), .Y(n917) );
  OAI22XL U1324 ( .A0(n523), .A1(n270), .B0(n1137), .B1(n1179), .Y(n918) );
  OAI22XL U1325 ( .A0(n524), .A1(n274), .B0(n1109), .B1(n1180), .Y(n919) );
  OAI22XL U1326 ( .A0(n525), .A1(n280), .B0(n1134), .B1(n1180), .Y(n920) );
  OAI22XL U1327 ( .A0(n526), .A1(n258), .B0(n1114), .B1(n1179), .Y(n921) );
  OAI22XL U1328 ( .A0(n527), .A1(n241), .B0(n1110), .B1(n1180), .Y(n922) );
  OAI22XL U1329 ( .A0(n528), .A1(n277), .B0(n1144), .B1(n1179), .Y(n923) );
  OAI22XL U1330 ( .A0(n529), .A1(n272), .B0(n1112), .B1(n1180), .Y(n924) );
  OAI22XL U1331 ( .A0(n530), .A1(n267), .B0(n1147), .B1(n1180), .Y(n925) );
  OAI22XL U1332 ( .A0(n531), .A1(n260), .B0(n1141), .B1(n1180), .Y(n926) );
  OAI22XL U1333 ( .A0(n532), .A1(n249), .B0(n1143), .B1(n1180), .Y(n927) );
  OAI22XL U1334 ( .A0(n533), .A1(n288), .B0(n1149), .B1(n1180), .Y(n928) );
  OAI22XL U1335 ( .A0(n534), .A1(n282), .B0(n1146), .B1(n1179), .Y(n929) );
  OAI22XL U1336 ( .A0(n535), .A1(n186), .B0(n1125), .B1(n1208), .Y(n931) );
  OAI22XL U1337 ( .A0(n536), .A1(n192), .B0(n1126), .B1(n1208), .Y(n932) );
  OAI22XL U1338 ( .A0(n537), .A1(n196), .B0(n1124), .B1(n1208), .Y(n933) );
  OAI22XL U1339 ( .A0(n538), .A1(n200), .B0(n1123), .B1(n1208), .Y(n934) );
  OAI22XL U1340 ( .A0(n539), .A1(n205), .B0(n1138), .B1(n1209), .Y(n935) );
  OAI22XL U1341 ( .A0(n540), .A1(n209), .B0(n1140), .B1(n1209), .Y(n936) );
  OAI22XL U1342 ( .A0(n541), .A1(n214), .B0(n1135), .B1(n1209), .Y(n937) );
  OAI22XL U1343 ( .A0(n542), .A1(n218), .B0(n1132), .B1(n1209), .Y(n938) );
  OAI22XL U1344 ( .A0(n543), .A1(n224), .B0(n1117), .B1(n1209), .Y(n939) );
  OAI22XL U1345 ( .A0(n544), .A1(n143), .B0(n1121), .B1(n1207), .Y(n940) );
  OAI22XL U1346 ( .A0(n545), .A1(n157), .B0(n1116), .B1(n1207), .Y(n941) );
  OAI22XL U1347 ( .A0(n546), .A1(n165), .B0(n1115), .B1(n1207), .Y(n942) );
  OAI22XL U1348 ( .A0(n547), .A1(n172), .B0(n1105), .B1(n1207), .Y(n943) );
  OAI22XL U1349 ( .A0(n548), .A1(n178), .B0(n1106), .B1(n1207), .Y(n944) );
  OAI22XL U1350 ( .A0(n549), .A1(n188), .B0(n1104), .B1(n1208), .Y(n945) );
  OAI22XL U1351 ( .A0(n550), .A1(n160), .B0(n1103), .B1(n1207), .Y(n946) );
  OAI22XL U1352 ( .A0(n551), .A1(n140), .B0(n1107), .B1(n146), .Y(n947) );
  OAI22XL U1353 ( .A0(n552), .A1(n181), .B0(n1108), .B1(n1208), .Y(n948) );
  OAI22XL U1354 ( .A0(n553), .A1(n175), .B0(n1113), .B1(n1207), .Y(n949) );
  OAI22XL U1355 ( .A0(n554), .A1(n168), .B0(n1111), .B1(n1207), .Y(n950) );
  OAI22XL U1356 ( .A0(n555), .A1(n162), .B0(n1122), .B1(n1207), .Y(n951) );
  OAI22XL U1357 ( .A0(n556), .A1(n148), .B0(n1118), .B1(n1207), .Y(n952) );
  OAI22XL U1358 ( .A0(n557), .A1(n227), .B0(n1120), .B1(n146), .Y(n953) );
  OAI22XL U1359 ( .A0(n558), .A1(n220), .B0(n1119), .B1(n1209), .Y(n954) );
  OAI22XL U1360 ( .A0(n559), .A1(n216), .B0(n1142), .B1(n1209), .Y(n955) );
  OAI22XL U1361 ( .A0(n560), .A1(n211), .B0(n1145), .B1(n1209), .Y(n956) );
  OAI22XL U1362 ( .A0(n561), .A1(n207), .B0(n1150), .B1(n1209), .Y(n957) );
  OAI22XL U1363 ( .A0(n562), .A1(n202), .B0(n1148), .B1(n1209), .Y(n958) );
  OAI22XL U1364 ( .A0(n563), .A1(n198), .B0(n1127), .B1(n1208), .Y(n959) );
  OAI22XL U1365 ( .A0(n564), .A1(n194), .B0(n1128), .B1(n1208), .Y(n960) );
  OAI22XL U1366 ( .A0(n565), .A1(n190), .B0(n1130), .B1(n1208), .Y(n961) );
  OAI22XL U1367 ( .A0(n566), .A1(n183), .B0(n1129), .B1(n1208), .Y(n962) );
  OAI22XL U1368 ( .A0(n567), .A1(n285), .B0(n1136), .B1(n1178), .Y(n963) );
  OAI22XL U1369 ( .A0(n568), .A1(n244), .B0(n1139), .B1(n1177), .Y(n964) );
  OAI22XL U1370 ( .A0(n569), .A1(n256), .B0(n1133), .B1(n1177), .Y(n965) );
  OAI22XL U1371 ( .A0(n570), .A1(n263), .B0(n1131), .B1(n1177), .Y(n966) );
  OAI22XL U1372 ( .A0(n571), .A1(n270), .B0(n1137), .B1(n1177), .Y(n967) );
  OAI22XL U1373 ( .A0(n572), .A1(n274), .B0(n1109), .B1(n1177), .Y(n968) );
  OAI22XL U1374 ( .A0(n573), .A1(n280), .B0(n1134), .B1(n1178), .Y(n969) );
  OAI22XL U1375 ( .A0(n574), .A1(n258), .B0(n1114), .B1(n1178), .Y(n970) );
  OAI22XL U1376 ( .A0(n575), .A1(n241), .B0(n1110), .B1(n1177), .Y(n971) );
  OAI22XL U1377 ( .A0(n576), .A1(n277), .B0(n1144), .B1(n1177), .Y(n972) );
  OAI22XL U1378 ( .A0(n577), .A1(n272), .B0(n1112), .B1(n1178), .Y(n973) );
  OAI22XL U1379 ( .A0(n578), .A1(n267), .B0(n1147), .B1(n1178), .Y(n974) );
  OAI22XL U1380 ( .A0(n579), .A1(n260), .B0(n1141), .B1(n1178), .Y(n975) );
  OAI22XL U1381 ( .A0(n580), .A1(n249), .B0(n1143), .B1(n1178), .Y(n976) );
  OAI22XL U1382 ( .A0(n581), .A1(n288), .B0(n1149), .B1(n1178), .Y(n977) );
  OAI22XL U1383 ( .A0(n582), .A1(n282), .B0(n1146), .B1(n1177), .Y(n978) );
  OAI22XL U1384 ( .A0(n584), .A1(n186), .B0(n1125), .B1(n1205), .Y(n981) );
  OAI22XL U1385 ( .A0(n585), .A1(n192), .B0(n1126), .B1(n1205), .Y(n982) );
  OAI22XL U1386 ( .A0(n586), .A1(n196), .B0(n1124), .B1(n1205), .Y(n983) );
  OAI22XL U1387 ( .A0(n587), .A1(n200), .B0(n1123), .B1(n1205), .Y(n984) );
  OAI22XL U1388 ( .A0(n588), .A1(n205), .B0(n1138), .B1(n1206), .Y(n985) );
  OAI22XL U1389 ( .A0(n589), .A1(n209), .B0(n1140), .B1(n1206), .Y(n986) );
  OAI22XL U1390 ( .A0(n590), .A1(n214), .B0(n1135), .B1(n1206), .Y(n987) );
  OAI22XL U1391 ( .A0(n591), .A1(n218), .B0(n1132), .B1(n1206), .Y(n988) );
  OAI22XL U1392 ( .A0(n592), .A1(n224), .B0(n1117), .B1(n1206), .Y(n989) );
  OAI22XL U1393 ( .A0(n593), .A1(n143), .B0(n1121), .B1(n1204), .Y(n990) );
  OAI22XL U1394 ( .A0(n594), .A1(n157), .B0(n1116), .B1(n1204), .Y(n991) );
  OAI22XL U1395 ( .A0(n595), .A1(n165), .B0(n1115), .B1(n1204), .Y(n992) );
  OAI22XL U1396 ( .A0(n596), .A1(n172), .B0(n1105), .B1(n1204), .Y(n993) );
  OAI22XL U1397 ( .A0(n597), .A1(n178), .B0(n1106), .B1(n1204), .Y(n994) );
  OAI22XL U1398 ( .A0(n598), .A1(n188), .B0(n1104), .B1(n1206), .Y(n995) );
  OAI22XL U1399 ( .A0(n599), .A1(n160), .B0(n1103), .B1(n147), .Y(n996) );
  OAI22XL U1400 ( .A0(n600), .A1(n140), .B0(n1107), .B1(n1204), .Y(n997) );
  OAI22XL U1401 ( .A0(n601), .A1(n181), .B0(n1108), .B1(n1205), .Y(n998) );
  OAI22XL U1402 ( .A0(n602), .A1(n175), .B0(n1113), .B1(n1204), .Y(n999) );
  OAI22XL U1403 ( .A0(n603), .A1(n168), .B0(n1111), .B1(n1204), .Y(n1000) );
  OAI22XL U1404 ( .A0(n604), .A1(n162), .B0(n1122), .B1(n1204), .Y(n1001) );
  OAI22XL U1405 ( .A0(n605), .A1(n148), .B0(n1118), .B1(n1204), .Y(n1002) );
  OAI22XL U1406 ( .A0(n606), .A1(n227), .B0(n1120), .B1(n147), .Y(n1003) );
  OAI22XL U1407 ( .A0(n607), .A1(n220), .B0(n1119), .B1(n1206), .Y(n1004) );
  OAI22XL U1408 ( .A0(n608), .A1(n216), .B0(n1142), .B1(n1206), .Y(n1005) );
  OAI22XL U1409 ( .A0(n609), .A1(n211), .B0(n1145), .B1(n1206), .Y(n1006) );
  OAI22XL U1410 ( .A0(n610), .A1(n207), .B0(n1150), .B1(n1206), .Y(n1007) );
  OAI22XL U1411 ( .A0(n611), .A1(n202), .B0(n1148), .B1(n1205), .Y(n1008) );
  OAI22XL U1412 ( .A0(n612), .A1(n198), .B0(n1127), .B1(n1205), .Y(n1009) );
  OAI22XL U1413 ( .A0(n613), .A1(n194), .B0(n1128), .B1(n1205), .Y(n1010) );
  OAI22XL U1414 ( .A0(n614), .A1(n190), .B0(n1130), .B1(n1205), .Y(n1011) );
  OAI22XL U1415 ( .A0(n615), .A1(n183), .B0(n1129), .B1(n1205), .Y(n1012) );
  OAI22XL U1416 ( .A0(n616), .A1(n285), .B0(n1136), .B1(n1165), .Y(n1013) );
  OAI22XL U1417 ( .A0(n617), .A1(n244), .B0(n1139), .B1(n1164), .Y(n1014) );
  OAI22XL U1418 ( .A0(n618), .A1(n256), .B0(n1133), .B1(n1165), .Y(n1015) );
  OAI22XL U1419 ( .A0(n619), .A1(n263), .B0(n1131), .B1(n1165), .Y(n1016) );
  OAI22XL U1420 ( .A0(n620), .A1(n270), .B0(n1137), .B1(n1165), .Y(n1017) );
  OAI22XL U1421 ( .A0(n621), .A1(n274), .B0(n1109), .B1(n1165), .Y(n1018) );
  OAI22XL U1422 ( .A0(n622), .A1(n280), .B0(n1134), .B1(n1165), .Y(n1019) );
  OAI22XL U1423 ( .A0(n623), .A1(n241), .B0(n1110), .B1(n1165), .Y(n1020) );
  OAI22XL U1424 ( .A0(n624), .A1(n277), .B0(n1144), .B1(n1164), .Y(n1021) );
  OAI22XL U1425 ( .A0(n625), .A1(n272), .B0(n1112), .B1(n1164), .Y(n1022) );
  OAI22XL U1426 ( .A0(n626), .A1(n267), .B0(n1147), .B1(n1164), .Y(n1023) );
  OAI22XL U1427 ( .A0(n627), .A1(n260), .B0(n1141), .B1(n1164), .Y(n1024) );
  OAI22XL U1428 ( .A0(n628), .A1(n249), .B0(n1143), .B1(n1164), .Y(n1025) );
  OAI22XL U1429 ( .A0(n629), .A1(n288), .B0(n1149), .B1(n1164), .Y(n1026) );
  OAI22XL U1430 ( .A0(n630), .A1(n282), .B0(n1146), .B1(n1164), .Y(n1027) );
  OAI22XL U1431 ( .A0(n631), .A1(n263), .B0(n1131), .B1(n1176), .Y(n1029) );
  OAI22XL U1432 ( .A0(n632), .A1(n258), .B0(n1114), .B1(n1176), .Y(n1030) );
  OAI22XL U1433 ( .A0(n633), .A1(n160), .B0(n1103), .B1(n1214), .Y(n1031) );
  OAI22XL U1434 ( .A0(n634), .A1(n165), .B0(n1115), .B1(n1213), .Y(n1032) );
  OAI22XL U1435 ( .A0(n635), .A1(n218), .B0(n1132), .B1(n1215), .Y(n1033) );
  OAI22XL U1436 ( .A0(n636), .A1(n200), .B0(n1123), .B1(n1214), .Y(n1034) );
  OAI22XL U1437 ( .A0(n637), .A1(n256), .B0(n1133), .B1(n1176), .Y(n1035) );
  OAI22XL U1438 ( .A0(n638), .A1(n280), .B0(n1134), .B1(n1175), .Y(n1036) );
  OAI22XL U1439 ( .A0(n639), .A1(n188), .B0(n1104), .B1(n1215), .Y(n1037) );
  OAI22XL U1440 ( .A0(n640), .A1(n157), .B0(n1116), .B1(n1213), .Y(n1038) );
  OAI22XL U1441 ( .A0(n641), .A1(n214), .B0(n1135), .B1(n1215), .Y(n1039) );
  OAI22XL U1442 ( .A0(n642), .A1(n196), .B0(n1124), .B1(n1214), .Y(n1040) );
  OAI22XL U1443 ( .A0(n643), .A1(n285), .B0(n1136), .B1(n1175), .Y(n1041) );
  OAI22XL U1444 ( .A0(n644), .A1(n270), .B0(n1137), .B1(n1176), .Y(n1042) );
  OAI22XL U1445 ( .A0(n645), .A1(n172), .B0(n1105), .B1(n1213), .Y(n1043) );
  OAI22XL U1446 ( .A0(n646), .A1(n224), .B0(n1117), .B1(n142), .Y(n1044) );
  OAI22XL U1447 ( .A0(n647), .A1(n205), .B0(n1138), .B1(n1215), .Y(n1045) );
  OAI22XL U1448 ( .A0(n648), .A1(n186), .B0(n1125), .B1(n1214), .Y(n1046) );
  OAI22XL U1449 ( .A0(n649), .A1(n244), .B0(n1139), .B1(n1176), .Y(n1047) );
  OAI22XL U1450 ( .A0(n650), .A1(n274), .B0(n1109), .B1(n1176), .Y(n1048) );
  OAI22XL U1451 ( .A0(n651), .A1(n178), .B0(n1106), .B1(n1213), .Y(n1049) );
  OAI22XL U1452 ( .A0(n652), .A1(n143), .B0(n1121), .B1(n1213), .Y(n1050) );
  OAI22XL U1453 ( .A0(n653), .A1(n209), .B0(n1140), .B1(n1215), .Y(n1051) );
  OAI22XL U1454 ( .A0(n654), .A1(n192), .B0(n1126), .B1(n1214), .Y(n1052) );
  OAI22XL U1455 ( .A0(n655), .A1(n260), .B0(n1141), .B1(n1175), .Y(n1053) );
  OAI22XL U1456 ( .A0(n656), .A1(n241), .B0(n1110), .B1(n1175), .Y(n1054) );
  OAI22XL U1457 ( .A0(n657), .A1(n140), .B0(n1107), .B1(n1213), .Y(n1055) );
  OAI22XL U1458 ( .A0(n658), .A1(n162), .B0(n1122), .B1(n1213), .Y(n1056) );
  OAI22XL U1459 ( .A0(n659), .A1(n216), .B0(n1142), .B1(n1215), .Y(n1057) );
  OAI22XL U1460 ( .A0(n660), .A1(n198), .B0(n1127), .B1(n1214), .Y(n1058) );
  OAI22XL U1461 ( .A0(n661), .A1(n249), .B0(n1143), .B1(n1175), .Y(n1059) );
  OAI22XL U1462 ( .A0(n662), .A1(n277), .B0(n1144), .B1(n1175), .Y(n1060) );
  OAI22XL U1463 ( .A0(n663), .A1(n181), .B0(n1108), .B1(n1214), .Y(n1061) );
  OAI22XL U1464 ( .A0(n664), .A1(n148), .B0(n1118), .B1(n1213), .Y(n1062) );
  OAI22XL U1465 ( .A0(n665), .A1(n211), .B0(n1145), .B1(n1215), .Y(n1063) );
  OAI22XL U1466 ( .A0(n666), .A1(n194), .B0(n1128), .B1(n1214), .Y(n1064) );
  OAI22XL U1467 ( .A0(n667), .A1(n282), .B0(n1146), .B1(n1176), .Y(n1065) );
  OAI22XL U1468 ( .A0(n668), .A1(n267), .B0(n1147), .B1(n1175), .Y(n1066) );
  OAI22XL U1469 ( .A0(n669), .A1(n168), .B0(n1111), .B1(n1213), .Y(n1067) );
  OAI22XL U1470 ( .A0(n670), .A1(n220), .B0(n1119), .B1(n1215), .Y(n1068) );
  OAI22XL U1471 ( .A0(n671), .A1(n202), .B0(n1148), .B1(n1215), .Y(n1069) );
  OAI22XL U1472 ( .A0(n672), .A1(n183), .B0(n1129), .B1(n1214), .Y(n1070) );
  OAI22XL U1473 ( .A0(n673), .A1(n288), .B0(n1149), .B1(n1176), .Y(n1071) );
  OAI22XL U1474 ( .A0(n674), .A1(n272), .B0(n1112), .B1(n1175), .Y(n1072) );
  OAI22XL U1475 ( .A0(n675), .A1(n175), .B0(n1113), .B1(n1213), .Y(n1073) );
  OAI22XL U1476 ( .A0(n676), .A1(n227), .B0(n1120), .B1(n142), .Y(n1074) );
  OAI22XL U1477 ( .A0(n677), .A1(n207), .B0(n1150), .B1(n1215), .Y(n1075) );
  OAI22XL U1478 ( .A0(n678), .A1(n190), .B0(n1130), .B1(n1214), .Y(n1076) );
  OAI22XL U1479 ( .A0(n685), .A1(n258), .B0(n1114), .B1(n1165), .Y(n1088) );
  OAI22XL U1480 ( .A0(n363), .A1(n162), .B0(n1122), .B1(n1198), .Y(n755) );
  OAI22XL U1481 ( .A0(n355), .A1(n172), .B0(n1105), .B1(n1198), .Y(n747) );
  NAND2X1 U1482 ( .A(n266), .B(n683), .Y(n255) );
  NAND2X1 U1483 ( .A(n276), .B(n683), .Y(n284) );
  NAND2X1 U1484 ( .A(data[7]), .B(n1182), .Y(n150) );
  NAND2X1 U1485 ( .A(data[6]), .B(n1183), .Y(n151) );
  NAND2X1 U1486 ( .A(data[5]), .B(n1183), .Y(n152) );
  NAND2X1 U1487 ( .A(data[4]), .B(n1183), .Y(n153) );
  NAND2X1 U1488 ( .A(data[3]), .B(n1182), .Y(n145) );
  NAND2X1 U1489 ( .A(data[2]), .B(n1182), .Y(n146) );
  NAND2X1 U1490 ( .A(data[0]), .B(n1183), .Y(n147) );
  NAND2X1 U1491 ( .A(data[1]), .B(n1182), .Y(n142) );
  NOR2X1 U1492 ( .A(n1181), .B(n680), .Y(n116) );
  NOR2X1 U1493 ( .A(n682), .B(n681), .Y(n29) );
  NOR2X1 U1494 ( .A(cnt_32[0]), .B(n681), .Y(n26) );
  OAI2BB2XL U1495 ( .B0(n683), .B1(n235), .A0N(N99), .A1N(n236), .Y(n1077) );
  NAND2X1 U1496 ( .A(phase[2]), .B(n233), .Y(n130) );
  OAI2BB2XL U1497 ( .B0(n680), .B1(n235), .A0N(N98), .A1N(n236), .Y(n1078) );
  OAI2BB2XL U1498 ( .B0(n682), .B1(n235), .A0N(n682), .A1N(n236), .Y(n1085) );
  OAI2BB2XL U1499 ( .B0(n684), .B1(n235), .A0N(N100), .A1N(n236), .Y(n1084) );
  OAI2BB2XL U1500 ( .B0(n681), .B1(n235), .A0N(N97), .A1N(n236), .Y(n1079) );
  OAI22XL U1501 ( .A0(n1320), .A1(n113), .B0(n1154), .B1(n121), .Y(n1083) );
  INVX1 U1502 ( .A(n121), .Y(n1320) );
  AND2X2 U1503 ( .A(n291), .B(n680), .Y(n276) );
  ADDHXL U1504 ( .A(cnt_32[1]), .B(cnt_32[0]), .CO(\r80/carry[2] ), .S(N97) );
  ADDHXL U1505 ( .A(cnt_32[2]), .B(\r80/carry[2] ), .CO(\r80/carry[3] ), .S(
        N98) );
  AND2X2 U1506 ( .A(n1323), .B(data[7]), .Y(n1155) );
  AND2X2 U1507 ( .A(n1323), .B(data[6]), .Y(n1156) );
  AND2X2 U1508 ( .A(n1323), .B(data[5]), .Y(n1157) );
  AND2X2 U1509 ( .A(n1323), .B(data[4]), .Y(n1158) );
  AND2X2 U1510 ( .A(n1323), .B(data[3]), .Y(n1159) );
  AND2X2 U1511 ( .A(n1323), .B(data[2]), .Y(n1160) );
  AND2X2 U1512 ( .A(n1323), .B(data[1]), .Y(n1161) );
  AND2X2 U1513 ( .A(n1323), .B(data[0]), .Y(n1162) );
  OAI32X1 U1514 ( .A0(n1324), .A1(n583), .A2(n137), .B0(n138), .B1(n1332), .Y(
        n980) );
  OAI32X1 U1515 ( .A0(n1324), .A1(n679), .A2(n137), .B0(n138), .B1(n1326), .Y(
        n1086) );
  OAI221XL U1516 ( .A0(result[23]), .A1(n18), .B0(result[55]), .B1(n19), .C0(
        n23), .Y(n15) );
  OA22X1 U1517 ( .A0(result[87]), .A1(n21), .B0(result[119]), .B1(n1218), .Y(
        n23) );
  OAI221XL U1518 ( .A0(result[22]), .A1(n1227), .B0(result[54]), .B1(n1224), 
        .C0(n37), .Y(n34) );
  OA22X1 U1519 ( .A0(result[86]), .A1(n1221), .B0(result[118]), .B1(n1217), 
        .Y(n37) );
  OAI221XL U1520 ( .A0(result[21]), .A1(n1226), .B0(result[53]), .B1(n1223), 
        .C0(n49), .Y(n46) );
  OA22X1 U1521 ( .A0(result[85]), .A1(n1220), .B0(result[117]), .B1(n22), .Y(
        n49) );
  OAI221XL U1522 ( .A0(result[20]), .A1(n1226), .B0(result[52]), .B1(n1223), 
        .C0(n61), .Y(n58) );
  OA22X1 U1523 ( .A0(result[84]), .A1(n1220), .B0(result[116]), .B1(n1218), 
        .Y(n61) );
  OAI221XL U1524 ( .A0(result[19]), .A1(n1227), .B0(result[51]), .B1(n1224), 
        .C0(n73), .Y(n70) );
  OA22X1 U1525 ( .A0(result[83]), .A1(n1221), .B0(result[115]), .B1(n1217), 
        .Y(n73) );
  OAI221XL U1526 ( .A0(result[18]), .A1(n1227), .B0(result[50]), .B1(n1224), 
        .C0(n85), .Y(n82) );
  OA22X1 U1527 ( .A0(result[82]), .A1(n1221), .B0(result[114]), .B1(n1217), 
        .Y(n85) );
  OAI221XL U1528 ( .A0(result[16]), .A1(n1227), .B0(result[48]), .B1(n1224), 
        .C0(n109), .Y(n106) );
  OA22X1 U1529 ( .A0(result[80]), .A1(n1221), .B0(result[112]), .B1(n1217), 
        .Y(n109) );
  OAI221XL U1530 ( .A0(result[17]), .A1(n1227), .B0(result[49]), .B1(n1224), 
        .C0(n97), .Y(n94) );
  OA22X1 U1531 ( .A0(result[81]), .A1(n1221), .B0(result[113]), .B1(n1217), 
        .Y(n97) );
  OAI221XL U1532 ( .A0(result[31]), .A1(n18), .B0(result[63]), .B1(n19), .C0(
        n20), .Y(n17) );
  OA22X1 U1533 ( .A0(result[95]), .A1(n21), .B0(result[127]), .B1(n1218), .Y(
        n20) );
  OAI221XL U1534 ( .A0(result[30]), .A1(n1227), .B0(result[62]), .B1(n1224), 
        .C0(n36), .Y(n35) );
  OA22X1 U1535 ( .A0(result[94]), .A1(n1221), .B0(result[126]), .B1(n1217), 
        .Y(n36) );
  OAI221XL U1536 ( .A0(result[29]), .A1(n1227), .B0(result[61]), .B1(n1224), 
        .C0(n48), .Y(n47) );
  OA22X1 U1537 ( .A0(result[93]), .A1(n1221), .B0(result[125]), .B1(n1217), 
        .Y(n48) );
  OAI221XL U1538 ( .A0(result[28]), .A1(n1226), .B0(result[60]), .B1(n1223), 
        .C0(n60), .Y(n59) );
  OA22X1 U1539 ( .A0(result[92]), .A1(n1220), .B0(result[124]), .B1(n22), .Y(
        n60) );
  OAI221XL U1540 ( .A0(result[27]), .A1(n1226), .B0(result[59]), .B1(n1223), 
        .C0(n72), .Y(n71) );
  OA22X1 U1541 ( .A0(result[91]), .A1(n1220), .B0(result[123]), .B1(n1218), 
        .Y(n72) );
  OAI221XL U1542 ( .A0(result[26]), .A1(n1227), .B0(result[58]), .B1(n1224), 
        .C0(n84), .Y(n83) );
  OA22X1 U1543 ( .A0(result[90]), .A1(n1221), .B0(result[122]), .B1(n1217), 
        .Y(n84) );
  OAI221XL U1544 ( .A0(result[24]), .A1(n1227), .B0(result[56]), .B1(n1224), 
        .C0(n108), .Y(n107) );
  OA22X1 U1545 ( .A0(result[88]), .A1(n1221), .B0(result[120]), .B1(n1217), 
        .Y(n108) );
  OAI221XL U1546 ( .A0(result[25]), .A1(n1227), .B0(result[57]), .B1(n1224), 
        .C0(n96), .Y(n95) );
  OA22X1 U1547 ( .A0(result[89]), .A1(n1221), .B0(result[121]), .B1(n1217), 
        .Y(n96) );
  ADDHXL U1548 ( .A(cnt_32[3]), .B(\r80/carry[3] ), .CO(\r80/carry[4] ), .S(
        N99) );
  XOR2X1 U1549 ( .A(\r80/carry[4] ), .B(cnt_32[4]), .Y(N100) );
  NAND4X1 U1550 ( .A(cnt_32[0]), .B(cnt_32[1]), .C(cnt_32[3]), .D(cnt_32[2]), 
        .Y(n1317) );
  NOR2BX1 U1551 ( .AN(n1317), .B(cnt_32[4]), .Y(N108) );
  AND4X1 U1552 ( .A(cnt_32[3]), .B(cnt_32[2]), .C(cnt_32[0]), .D(cnt_32[1]), 
        .Y(n1319) );
  OAI21XL U1553 ( .A0(cnt_32[4]), .A1(n1319), .B0(n1318), .Y(N94) );
endmodule

